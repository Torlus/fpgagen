-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM1;

architecture arch of CtrlROM_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"ac080b0b",
    10 => x"0bbdb008",
    11 => x"0b0b0bbd",
    12 => x"b4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bdb40c0b",
    16 => x"0b0bbdb0",
    17 => x"0c0b0b0b",
    18 => x"bdac0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb7b0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bdac7080",
    57 => x"c7ec278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518f9a04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbdbc0c",
    65 => x"9f0bbdc0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bdc008ff",
    69 => x"05bdc00c",
    70 => x"bdc00880",
    71 => x"25eb38bd",
    72 => x"bc08ff05",
    73 => x"bdbc0cbd",
    74 => x"bc088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbd",
    94 => x"bc08258f",
    95 => x"3882b32d",
    96 => x"bdbc08ff",
    97 => x"05bdbc0c",
    98 => x"82f504bd",
    99 => x"bc08bdc0",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038bdbc",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"bdc00881",
   109 => x"05bdc00c",
   110 => x"bdc00851",
   111 => x"9f7125e2",
   112 => x"38800bbd",
   113 => x"c00cbdbc",
   114 => x"088105bd",
   115 => x"bc0c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34bdc008",
   120 => x"8105bdc0",
   121 => x"0cbdc008",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbdc00c",
   125 => x"bdbc0881",
   126 => x"05bdbc0c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"bdc40cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbd",
   162 => x"c40c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72bdc408",
   167 => x"8407bdc4",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"baac0c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"bdc40852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c7d00cba",
   200 => x"cc718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"bdac0c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b8c452bd",
   211 => x"c8519c8d",
   212 => x"2dbdac08",
   213 => x"802ea138",
   214 => x"80c0e452",
   215 => x"bdc8519e",
   216 => x"ce2d80c0",
   217 => x"e408bdd4",
   218 => x"0c80c0e4",
   219 => x"08fec00c",
   220 => x"80c0e408",
   221 => x"5186932d",
   222 => x"0288050d",
   223 => x"0402f005",
   224 => x"0d805191",
   225 => x"dc2db8c4",
   226 => x"52bdc851",
   227 => x"9c8d2dbd",
   228 => x"ac08802e",
   229 => x"a838bdd4",
   230 => x"0880c0e4",
   231 => x"0c80c0e8",
   232 => x"5480fd53",
   233 => x"80747084",
   234 => x"05560cff",
   235 => x"13537280",
   236 => x"25f23880",
   237 => x"c0e452bd",
   238 => x"c8519ef7",
   239 => x"2d029005",
   240 => x"0d0402d8",
   241 => x"050d800b",
   242 => x"bab00cbd",
   243 => x"d408fec0",
   244 => x"0c810bfe",
   245 => x"c40c840b",
   246 => x"fec40c7b",
   247 => x"52bdc851",
   248 => x"9c8d2dbd",
   249 => x"ac0853bd",
   250 => x"ac08802e",
   251 => x"81b338bd",
   252 => x"cc085580",
   253 => x"0bff1657",
   254 => x"5975792e",
   255 => x"8b388119",
   256 => x"76812a57",
   257 => x"5975f738",
   258 => x"f7195974",
   259 => x"b080802e",
   260 => x"09810689",
   261 => x"38820bfe",
   262 => x"dc0c88b4",
   263 => x"04749880",
   264 => x"802e0981",
   265 => x"06893881",
   266 => x"0bfedc0c",
   267 => x"88b40480",
   268 => x"0bfedc0c",
   269 => x"815a8075",
   270 => x"2580df38",
   271 => x"78527551",
   272 => x"84812d80",
   273 => x"c0e452bd",
   274 => x"c8519ece",
   275 => x"2dbdac08",
   276 => x"802ea838",
   277 => x"80c0e458",
   278 => x"83fc5777",
   279 => x"70840559",
   280 => x"087083ff",
   281 => x"ff067190",
   282 => x"2afec80c",
   283 => x"fec80cfc",
   284 => x"18585376",
   285 => x"8025e438",
   286 => x"898204bd",
   287 => x"ac085a84",
   288 => x"8055bdc8",
   289 => x"519ea02d",
   290 => x"fc801581",
   291 => x"17575574",
   292 => x"8024ffa8",
   293 => x"3879802e",
   294 => x"8638820b",
   295 => x"bab00c79",
   296 => x"5372bdac",
   297 => x"0c02a805",
   298 => x"0d0402fc",
   299 => x"050dabf4",
   300 => x"2dfec451",
   301 => x"81710c82",
   302 => x"710c0284",
   303 => x"050d0402",
   304 => x"f4050d74",
   305 => x"76785354",
   306 => x"52807125",
   307 => x"97387270",
   308 => x"81055480",
   309 => x"f52d7270",
   310 => x"81055481",
   311 => x"b72dff11",
   312 => x"5170eb38",
   313 => x"807281b7",
   314 => x"2d028c05",
   315 => x"0d0402e8",
   316 => x"050d7756",
   317 => x"80705654",
   318 => x"737624b3",
   319 => x"3880c6f4",
   320 => x"08742eab",
   321 => x"38735199",
   322 => x"d62dbdac",
   323 => x"08bdac08",
   324 => x"09810570",
   325 => x"bdac0807",
   326 => x"9f2a7705",
   327 => x"81175757",
   328 => x"53537476",
   329 => x"24893880",
   330 => x"c6f40874",
   331 => x"26d73872",
   332 => x"bdac0c02",
   333 => x"98050d04",
   334 => x"02f4050d",
   335 => x"bcd80815",
   336 => x"5189ee2d",
   337 => x"bdac0880",
   338 => x"2e95388b",
   339 => x"53bdac08",
   340 => x"5280c4e4",
   341 => x"5189bf2d",
   342 => x"80c4e451",
   343 => x"87c22dba",
   344 => x"b451add8",
   345 => x"2dabf42d",
   346 => x"805184e6",
   347 => x"2d028c05",
   348 => x"0d0402dc",
   349 => x"050d8070",
   350 => x"5a5574bc",
   351 => x"d80825b1",
   352 => x"3880c6f4",
   353 => x"08752ea9",
   354 => x"38785199",
   355 => x"d62dbdac",
   356 => x"08098105",
   357 => x"70bdac08",
   358 => x"079f2a76",
   359 => x"05811b5b",
   360 => x"565474bc",
   361 => x"d8082589",
   362 => x"3880c6f4",
   363 => x"087926d9",
   364 => x"38805578",
   365 => x"80c6f408",
   366 => x"2781d038",
   367 => x"785199d6",
   368 => x"2dbdac08",
   369 => x"802e81a5",
   370 => x"38bdac08",
   371 => x"8b0580f5",
   372 => x"2d70842a",
   373 => x"70810677",
   374 => x"1078842b",
   375 => x"80c4e40b",
   376 => x"80f52d5c",
   377 => x"5c535155",
   378 => x"5673802e",
   379 => x"80c73874",
   380 => x"16822b8d",
   381 => x"ae0bbbac",
   382 => x"120c5477",
   383 => x"753110bd",
   384 => x"dc115556",
   385 => x"90747081",
   386 => x"055681b7",
   387 => x"2da07481",
   388 => x"b72d7681",
   389 => x"ff068116",
   390 => x"58547380",
   391 => x"2e8a389c",
   392 => x"5380c4e4",
   393 => x"528cae04",
   394 => x"8b53bdac",
   395 => x"0852bdde",
   396 => x"16518ce5",
   397 => x"04741682",
   398 => x"2b8ab80b",
   399 => x"bbac120c",
   400 => x"547681ff",
   401 => x"06811658",
   402 => x"5473802e",
   403 => x"8a389c53",
   404 => x"80c4e452",
   405 => x"8cdd048b",
   406 => x"53bdac08",
   407 => x"52777531",
   408 => x"10bddc05",
   409 => x"51765589",
   410 => x"bf2d8d80",
   411 => x"04749029",
   412 => x"75317010",
   413 => x"bddc0551",
   414 => x"54bdac08",
   415 => x"7481b72d",
   416 => x"81195974",
   417 => x"8b24a238",
   418 => x"8bb30474",
   419 => x"90297531",
   420 => x"7010bddc",
   421 => x"058c7731",
   422 => x"57515480",
   423 => x"7481b72d",
   424 => x"9e14ff16",
   425 => x"565474f3",
   426 => x"3802a405",
   427 => x"0d0402fc",
   428 => x"050dbcd8",
   429 => x"08135189",
   430 => x"ee2dbdac",
   431 => x"08802e88",
   432 => x"38bdac08",
   433 => x"5191dc2d",
   434 => x"800bbcd8",
   435 => x"0c8af22d",
   436 => x"acb72d02",
   437 => x"84050d04",
   438 => x"02fc050d",
   439 => x"725170fd",
   440 => x"2ead3870",
   441 => x"fd248a38",
   442 => x"70fc2e80",
   443 => x"c4388eb9",
   444 => x"0470fe2e",
   445 => x"b13870ff",
   446 => x"2e098106",
   447 => x"bc38bcd8",
   448 => x"08517080",
   449 => x"2eb338ff",
   450 => x"11bcd80c",
   451 => x"8eb904bc",
   452 => x"d808f005",
   453 => x"70bcd80c",
   454 => x"51708025",
   455 => x"9c38800b",
   456 => x"bcd80c8e",
   457 => x"b904bcd8",
   458 => x"088105bc",
   459 => x"d80c8eb9",
   460 => x"04bcd808",
   461 => x"9005bcd8",
   462 => x"0c8af22d",
   463 => x"acb72d02",
   464 => x"84050d04",
   465 => x"02fc050d",
   466 => x"800bbcd8",
   467 => x"0c8af22d",
   468 => x"bba451ad",
   469 => x"d82d0284",
   470 => x"050d0402",
   471 => x"f8050d80",
   472 => x"c7d00882",
   473 => x"06bad40b",
   474 => x"80f52d52",
   475 => x"5270802e",
   476 => x"85387181",
   477 => x"0752baec",
   478 => x"0b80f52d",
   479 => x"5170802e",
   480 => x"85387184",
   481 => x"0752bdd8",
   482 => x"08802e85",
   483 => x"38719007",
   484 => x"5271bdac",
   485 => x"0c028805",
   486 => x"0d0402f4",
   487 => x"050d810b",
   488 => x"bdd80c80",
   489 => x"0bbab00c",
   490 => x"90518693",
   491 => x"2d810bfe",
   492 => x"c40c840b",
   493 => x"fec40c83",
   494 => x"0bfecc0c",
   495 => x"b8d05185",
   496 => x"f22d8452",
   497 => x"a3ae2d92",
   498 => x"fd2dbdac",
   499 => x"08802e86",
   500 => x"38fe528f",
   501 => x"de04ff12",
   502 => x"52718024",
   503 => x"e7387180",
   504 => x"2e81ab38",
   505 => x"a9c02dab",
   506 => x"d52da9a3",
   507 => x"2da9a32d",
   508 => x"81f82d81",
   509 => x"5184e62d",
   510 => x"a9a32da9",
   511 => x"a32d8151",
   512 => x"84e62d86",
   513 => x"c42db8e8",
   514 => x"5187c22d",
   515 => x"bdac0880",
   516 => x"2e9438ba",
   517 => x"b451add8",
   518 => x"2d805184",
   519 => x"e62d820b",
   520 => x"bab00c90",
   521 => x"b004bdac",
   522 => x"08518ec4",
   523 => x"2dabe12d",
   524 => x"a9d92dad",
   525 => x"eb2dbdac",
   526 => x"0880c7d4",
   527 => x"08882b80",
   528 => x"c7d80807",
   529 => x"fed80c53",
   530 => x"8edb2dbd",
   531 => x"ac08bdd4",
   532 => x"082ea238",
   533 => x"bdac08bd",
   534 => x"d40cbdac",
   535 => x"08fec00c",
   536 => x"84527251",
   537 => x"84e62da9",
   538 => x"a32da9a3",
   539 => x"2dff1252",
   540 => x"718025ee",
   541 => x"3872802e",
   542 => x"8c38bab0",
   543 => x"088807fe",
   544 => x"c40c90b0",
   545 => x"04bab008",
   546 => x"fec40c90",
   547 => x"b004b8f4",
   548 => x"5185f22d",
   549 => x"800bbdac",
   550 => x"0c028c05",
   551 => x"0d0402e8",
   552 => x"050d7779",
   553 => x"7b585555",
   554 => x"80537276",
   555 => x"25a33874",
   556 => x"70810556",
   557 => x"80f52d74",
   558 => x"70810556",
   559 => x"80f52d52",
   560 => x"5271712e",
   561 => x"86388151",
   562 => x"91d30481",
   563 => x"135391aa",
   564 => x"04805170",
   565 => x"bdac0c02",
   566 => x"98050d04",
   567 => x"02ec050d",
   568 => x"76557480",
   569 => x"2ebe389a",
   570 => x"1580e02d",
   571 => x"51a7e82d",
   572 => x"bdac08bd",
   573 => x"ac0880c7",
   574 => x"940cbdac",
   575 => x"08545480",
   576 => x"c6f00880",
   577 => x"2e993894",
   578 => x"1580e02d",
   579 => x"51a7e82d",
   580 => x"bdac0890",
   581 => x"2b83fff0",
   582 => x"0a067075",
   583 => x"07515372",
   584 => x"80c7940c",
   585 => x"80c79408",
   586 => x"5372802e",
   587 => x"9d3880c6",
   588 => x"e808fe14",
   589 => x"712980c6",
   590 => x"fc080580",
   591 => x"c7980c70",
   592 => x"842b80c6",
   593 => x"f40c5492",
   594 => x"f80480c7",
   595 => x"800880c7",
   596 => x"940c80c7",
   597 => x"840880c7",
   598 => x"980c80c6",
   599 => x"f008802e",
   600 => x"8b3880c6",
   601 => x"e808842b",
   602 => x"5392f304",
   603 => x"80c78808",
   604 => x"842b5372",
   605 => x"80c6f40c",
   606 => x"0294050d",
   607 => x"0402d805",
   608 => x"0d800b80",
   609 => x"c6f00c80",
   610 => x"c0e45280",
   611 => x"51a6982d",
   612 => x"bdac0854",
   613 => x"bdac088c",
   614 => x"38b98851",
   615 => x"85f22d73",
   616 => x"5598d904",
   617 => x"8056810b",
   618 => x"80c79c0c",
   619 => x"8853b994",
   620 => x"5280c19a",
   621 => x"51919e2d",
   622 => x"bdac0876",
   623 => x"2e098106",
   624 => x"8838bdac",
   625 => x"0880c79c",
   626 => x"0c8853b9",
   627 => x"a05280c1",
   628 => x"b651919e",
   629 => x"2dbdac08",
   630 => x"8838bdac",
   631 => x"0880c79c",
   632 => x"0c80c79c",
   633 => x"08802e80",
   634 => x"fd3880c4",
   635 => x"aa0b80f5",
   636 => x"2d80c4ab",
   637 => x"0b80f52d",
   638 => x"71982b71",
   639 => x"902b0780",
   640 => x"c4ac0b80",
   641 => x"f52d7088",
   642 => x"2b720780",
   643 => x"c4ad0b80",
   644 => x"f52d7107",
   645 => x"80c4e20b",
   646 => x"80f52d80",
   647 => x"c4e30b80",
   648 => x"f52d7188",
   649 => x"2b07535f",
   650 => x"54525a56",
   651 => x"57557381",
   652 => x"abaa2e09",
   653 => x"81068d38",
   654 => x"7551a7b8",
   655 => x"2dbdac08",
   656 => x"5694d104",
   657 => x"7382d4d5",
   658 => x"2e8738b9",
   659 => x"ac519596",
   660 => x"0480c0e4",
   661 => x"527551a6",
   662 => x"982dbdac",
   663 => x"0855bdac",
   664 => x"08802e83",
   665 => x"f4388853",
   666 => x"b9a05280",
   667 => x"c1b65191",
   668 => x"9e2dbdac",
   669 => x"088a3881",
   670 => x"0b80c6f0",
   671 => x"0c959c04",
   672 => x"8853b994",
   673 => x"5280c19a",
   674 => x"51919e2d",
   675 => x"bdac0880",
   676 => x"2e8a38b9",
   677 => x"c05185f2",
   678 => x"2d95fb04",
   679 => x"80c4e20b",
   680 => x"80f52d54",
   681 => x"7380d52e",
   682 => x"09810680",
   683 => x"ce3880c4",
   684 => x"e30b80f5",
   685 => x"2d547381",
   686 => x"aa2e0981",
   687 => x"06bd3880",
   688 => x"0b80c0e4",
   689 => x"0b80f52d",
   690 => x"56547481",
   691 => x"e92e8338",
   692 => x"81547481",
   693 => x"eb2e8c38",
   694 => x"80557375",
   695 => x"2e098106",
   696 => x"82f73880",
   697 => x"c0ef0b80",
   698 => x"f52d5574",
   699 => x"8e3880c0",
   700 => x"f00b80f5",
   701 => x"2d547382",
   702 => x"2e863880",
   703 => x"5598d904",
   704 => x"80c0f10b",
   705 => x"80f52d70",
   706 => x"80c6e80c",
   707 => x"ff0580c6",
   708 => x"ec0c80c0",
   709 => x"f20b80f5",
   710 => x"2d80c0f3",
   711 => x"0b80f52d",
   712 => x"58760577",
   713 => x"82802905",
   714 => x"7080c6f8",
   715 => x"0c80c0f4",
   716 => x"0b80f52d",
   717 => x"7080c78c",
   718 => x"0c80c6f0",
   719 => x"08595758",
   720 => x"76802e81",
   721 => x"b5388853",
   722 => x"b9a05280",
   723 => x"c1b65191",
   724 => x"9e2dbdac",
   725 => x"08828238",
   726 => x"80c6e808",
   727 => x"70842b80",
   728 => x"c6f40c70",
   729 => x"80c7880c",
   730 => x"80c1890b",
   731 => x"80f52d80",
   732 => x"c1880b80",
   733 => x"f52d7182",
   734 => x"80290580",
   735 => x"c18a0b80",
   736 => x"f52d7084",
   737 => x"80802912",
   738 => x"80c18b0b",
   739 => x"80f52d70",
   740 => x"81800a29",
   741 => x"127080c7",
   742 => x"900c80c7",
   743 => x"8c087129",
   744 => x"80c6f808",
   745 => x"057080c6",
   746 => x"fc0c80c1",
   747 => x"910b80f5",
   748 => x"2d80c190",
   749 => x"0b80f52d",
   750 => x"71828029",
   751 => x"0580c192",
   752 => x"0b80f52d",
   753 => x"70848080",
   754 => x"291280c1",
   755 => x"930b80f5",
   756 => x"2d70982b",
   757 => x"81f00a06",
   758 => x"72057080",
   759 => x"c7800cfe",
   760 => x"117e2977",
   761 => x"0580c784",
   762 => x"0c525952",
   763 => x"43545e51",
   764 => x"5259525d",
   765 => x"57595798",
   766 => x"d20480c0",
   767 => x"f60b80f5",
   768 => x"2d80c0f5",
   769 => x"0b80f52d",
   770 => x"71828029",
   771 => x"057080c6",
   772 => x"f40c70a0",
   773 => x"2983ff05",
   774 => x"70892a70",
   775 => x"80c7880c",
   776 => x"80c0fb0b",
   777 => x"80f52d80",
   778 => x"c0fa0b80",
   779 => x"f52d7182",
   780 => x"80290570",
   781 => x"80c7900c",
   782 => x"7b71291e",
   783 => x"7080c784",
   784 => x"0c7d80c7",
   785 => x"800c7305",
   786 => x"80c6fc0c",
   787 => x"555e5151",
   788 => x"55558051",
   789 => x"91dc2d81",
   790 => x"5574bdac",
   791 => x"0c02a805",
   792 => x"0d0402ec",
   793 => x"050d7670",
   794 => x"872c7180",
   795 => x"ff065556",
   796 => x"5480c6f0",
   797 => x"088a3873",
   798 => x"882c7481",
   799 => x"ff065455",
   800 => x"80c0e452",
   801 => x"80c6f808",
   802 => x"1551a698",
   803 => x"2dbdac08",
   804 => x"54bdac08",
   805 => x"802eb638",
   806 => x"80c6f008",
   807 => x"802e9938",
   808 => x"72842980",
   809 => x"c0e40570",
   810 => x"085253a7",
   811 => x"b82dbdac",
   812 => x"08f00a06",
   813 => x"5399cb04",
   814 => x"721080c0",
   815 => x"e4057080",
   816 => x"e02d5253",
   817 => x"a7e82dbd",
   818 => x"ac085372",
   819 => x"5473bdac",
   820 => x"0c029405",
   821 => x"0d0402e0",
   822 => x"050d7970",
   823 => x"842c80c7",
   824 => x"98080571",
   825 => x"8f065255",
   826 => x"53728a38",
   827 => x"80c0e452",
   828 => x"7351a698",
   829 => x"2d72a029",
   830 => x"80c0e405",
   831 => x"54807480",
   832 => x"f52d5653",
   833 => x"74732e83",
   834 => x"38815374",
   835 => x"81e52e81",
   836 => x"f1388170",
   837 => x"74065458",
   838 => x"72802e81",
   839 => x"e5388b14",
   840 => x"80f52d70",
   841 => x"832a7906",
   842 => x"58567699",
   843 => x"38bcdc08",
   844 => x"53728938",
   845 => x"7280c4e4",
   846 => x"0b81b72d",
   847 => x"76bcdc0c",
   848 => x"73539c84",
   849 => x"04758f2e",
   850 => x"09810681",
   851 => x"b538749f",
   852 => x"068d2980",
   853 => x"c4d71151",
   854 => x"53811480",
   855 => x"f52d7370",
   856 => x"81055581",
   857 => x"b72d8314",
   858 => x"80f52d73",
   859 => x"70810555",
   860 => x"81b72d85",
   861 => x"1480f52d",
   862 => x"73708105",
   863 => x"5581b72d",
   864 => x"871480f5",
   865 => x"2d737081",
   866 => x"055581b7",
   867 => x"2d891480",
   868 => x"f52d7370",
   869 => x"81055581",
   870 => x"b72d8e14",
   871 => x"80f52d73",
   872 => x"70810555",
   873 => x"81b72d90",
   874 => x"1480f52d",
   875 => x"73708105",
   876 => x"5581b72d",
   877 => x"921480f5",
   878 => x"2d737081",
   879 => x"055581b7",
   880 => x"2d941480",
   881 => x"f52d7370",
   882 => x"81055581",
   883 => x"b72d9614",
   884 => x"80f52d73",
   885 => x"70810555",
   886 => x"81b72d98",
   887 => x"1480f52d",
   888 => x"73708105",
   889 => x"5581b72d",
   890 => x"9c1480f5",
   891 => x"2d737081",
   892 => x"055581b7",
   893 => x"2d9e1480",
   894 => x"f52d7381",
   895 => x"b72d77bc",
   896 => x"dc0c8053",
   897 => x"72bdac0c",
   898 => x"02a0050d",
   899 => x"0402cc05",
   900 => x"0d7e605e",
   901 => x"5a800b80",
   902 => x"c7940880",
   903 => x"c7980859",
   904 => x"5c568058",
   905 => x"80c6f408",
   906 => x"782e81b2",
   907 => x"38778f06",
   908 => x"a0175754",
   909 => x"73913880",
   910 => x"c0e45276",
   911 => x"51811757",
   912 => x"a6982d80",
   913 => x"c0e45680",
   914 => x"7680f52d",
   915 => x"56547474",
   916 => x"2e833881",
   917 => x"547481e5",
   918 => x"2e80f738",
   919 => x"81707506",
   920 => x"555c7380",
   921 => x"2e80eb38",
   922 => x"8b1680f5",
   923 => x"2d980659",
   924 => x"7880df38",
   925 => x"8b537c52",
   926 => x"7551919e",
   927 => x"2dbdac08",
   928 => x"80d0389c",
   929 => x"160851a7",
   930 => x"b82dbdac",
   931 => x"08841b0c",
   932 => x"9a1680e0",
   933 => x"2d51a7e8",
   934 => x"2dbdac08",
   935 => x"bdac0888",
   936 => x"1c0cbdac",
   937 => x"08555580",
   938 => x"c6f00880",
   939 => x"2e983894",
   940 => x"1680e02d",
   941 => x"51a7e82d",
   942 => x"bdac0890",
   943 => x"2b83fff0",
   944 => x"0a067016",
   945 => x"51547388",
   946 => x"1b0c787a",
   947 => x"0c7b549e",
   948 => x"97048118",
   949 => x"5880c6f4",
   950 => x"087826fe",
   951 => x"d03880c6",
   952 => x"f008802e",
   953 => x"b0387a51",
   954 => x"98e22dbd",
   955 => x"ac08bdac",
   956 => x"0880ffff",
   957 => x"fff80655",
   958 => x"5b7380ff",
   959 => x"fffff82e",
   960 => x"9438bdac",
   961 => x"08fe0580",
   962 => x"c6e80829",
   963 => x"80c6fc08",
   964 => x"05579ca2",
   965 => x"04805473",
   966 => x"bdac0c02",
   967 => x"b4050d04",
   968 => x"02f4050d",
   969 => x"74700881",
   970 => x"05710c70",
   971 => x"0880c6ec",
   972 => x"08065353",
   973 => x"718e3888",
   974 => x"13085198",
   975 => x"e22dbdac",
   976 => x"0888140c",
   977 => x"810bbdac",
   978 => x"0c028c05",
   979 => x"0d0402f0",
   980 => x"050d7588",
   981 => x"1108fe05",
   982 => x"80c6e808",
   983 => x"2980c6fc",
   984 => x"08117208",
   985 => x"80c6ec08",
   986 => x"06057955",
   987 => x"535454a6",
   988 => x"982d0290",
   989 => x"050d0402",
   990 => x"f0050d75",
   991 => x"881108fe",
   992 => x"0580c6e8",
   993 => x"082980c6",
   994 => x"fc081172",
   995 => x"0880c6ec",
   996 => x"08060579",
   997 => x"55535454",
   998 => x"a4d82d02",
   999 => x"90050d04",
  1000 => x"02f4050d",
  1001 => x"d45281ff",
  1002 => x"720c7108",
  1003 => x"5381ff72",
  1004 => x"0c72882b",
  1005 => x"83fe8006",
  1006 => x"72087081",
  1007 => x"ff065152",
  1008 => x"5381ff72",
  1009 => x"0c727107",
  1010 => x"882b7208",
  1011 => x"7081ff06",
  1012 => x"51525381",
  1013 => x"ff720c72",
  1014 => x"7107882b",
  1015 => x"72087081",
  1016 => x"ff067207",
  1017 => x"bdac0c52",
  1018 => x"53028c05",
  1019 => x"0d0402f4",
  1020 => x"050d7476",
  1021 => x"7181ff06",
  1022 => x"d40c5353",
  1023 => x"80c7a008",
  1024 => x"85387189",
  1025 => x"2b527198",
  1026 => x"2ad40c71",
  1027 => x"902a7081",
  1028 => x"ff06d40c",
  1029 => x"5171882a",
  1030 => x"7081ff06",
  1031 => x"d40c5171",
  1032 => x"81ff06d4",
  1033 => x"0c72902a",
  1034 => x"7081ff06",
  1035 => x"d40c51d4",
  1036 => x"087081ff",
  1037 => x"06515182",
  1038 => x"b8bf5270",
  1039 => x"81ff2e09",
  1040 => x"81069438",
  1041 => x"81ff0bd4",
  1042 => x"0cd40870",
  1043 => x"81ff06ff",
  1044 => x"14545151",
  1045 => x"71e53870",
  1046 => x"bdac0c02",
  1047 => x"8c050d04",
  1048 => x"02fc050d",
  1049 => x"81c75181",
  1050 => x"ff0bd40c",
  1051 => x"ff115170",
  1052 => x"8025f438",
  1053 => x"0284050d",
  1054 => x"0402f005",
  1055 => x"0da0e02d",
  1056 => x"8fcf5380",
  1057 => x"5287fc80",
  1058 => x"f7519fee",
  1059 => x"2dbdac08",
  1060 => x"54bdac08",
  1061 => x"812e0981",
  1062 => x"06a33881",
  1063 => x"ff0bd40c",
  1064 => x"820a5284",
  1065 => x"9c80e951",
  1066 => x"9fee2dbd",
  1067 => x"ac088b38",
  1068 => x"81ff0bd4",
  1069 => x"0c7353a1",
  1070 => x"c304a0e0",
  1071 => x"2dff1353",
  1072 => x"72c13872",
  1073 => x"bdac0c02",
  1074 => x"90050d04",
  1075 => x"02f4050d",
  1076 => x"81ff0bd4",
  1077 => x"0c935380",
  1078 => x"5287fc80",
  1079 => x"c1519fee",
  1080 => x"2dbdac08",
  1081 => x"8b3881ff",
  1082 => x"0bd40c81",
  1083 => x"53a1f904",
  1084 => x"a0e02dff",
  1085 => x"135372df",
  1086 => x"3872bdac",
  1087 => x"0c028c05",
  1088 => x"0d0402f0",
  1089 => x"050da0e0",
  1090 => x"2d83aa52",
  1091 => x"849c80c8",
  1092 => x"519fee2d",
  1093 => x"bdac0881",
  1094 => x"2e098106",
  1095 => x"92389fa0",
  1096 => x"2dbdac08",
  1097 => x"83ffff06",
  1098 => x"537283aa",
  1099 => x"2e9738a1",
  1100 => x"cc2da2c0",
  1101 => x"048154a3",
  1102 => x"a504b9cc",
  1103 => x"5185f22d",
  1104 => x"8054a3a5",
  1105 => x"0481ff0b",
  1106 => x"d40cb153",
  1107 => x"a0f92dbd",
  1108 => x"ac08802e",
  1109 => x"80c03880",
  1110 => x"5287fc80",
  1111 => x"fa519fee",
  1112 => x"2dbdac08",
  1113 => x"b13881ff",
  1114 => x"0bd40cd4",
  1115 => x"085381ff",
  1116 => x"0bd40c81",
  1117 => x"ff0bd40c",
  1118 => x"81ff0bd4",
  1119 => x"0c81ff0b",
  1120 => x"d40c7286",
  1121 => x"2a708106",
  1122 => x"bdac0856",
  1123 => x"51537280",
  1124 => x"2e9338a2",
  1125 => x"b5047282",
  1126 => x"2eff9f38",
  1127 => x"ff135372",
  1128 => x"ffaa3872",
  1129 => x"5473bdac",
  1130 => x"0c029005",
  1131 => x"0d0402f0",
  1132 => x"050d810b",
  1133 => x"80c7a00c",
  1134 => x"8454d008",
  1135 => x"708f2a70",
  1136 => x"81065151",
  1137 => x"5372f338",
  1138 => x"72d00ca0",
  1139 => x"e02db9dc",
  1140 => x"5185f22d",
  1141 => x"d008708f",
  1142 => x"2a708106",
  1143 => x"51515372",
  1144 => x"f338810b",
  1145 => x"d00cb153",
  1146 => x"805284d4",
  1147 => x"80c0519f",
  1148 => x"ee2dbdac",
  1149 => x"08812ea1",
  1150 => x"3872822e",
  1151 => x"0981068c",
  1152 => x"38b9e851",
  1153 => x"85f22d80",
  1154 => x"53a4cf04",
  1155 => x"ff135372",
  1156 => x"d738ff14",
  1157 => x"5473ffa2",
  1158 => x"38a2822d",
  1159 => x"bdac0880",
  1160 => x"c7a00cbd",
  1161 => x"ac088b38",
  1162 => x"815287fc",
  1163 => x"80d0519f",
  1164 => x"ee2d81ff",
  1165 => x"0bd40cd0",
  1166 => x"08708f2a",
  1167 => x"70810651",
  1168 => x"515372f3",
  1169 => x"3872d00c",
  1170 => x"81ff0bd4",
  1171 => x"0c815372",
  1172 => x"bdac0c02",
  1173 => x"90050d04",
  1174 => x"02e8050d",
  1175 => x"785681ff",
  1176 => x"0bd40cd0",
  1177 => x"08708f2a",
  1178 => x"70810651",
  1179 => x"515372f3",
  1180 => x"3882810b",
  1181 => x"d00c81ff",
  1182 => x"0bd40c77",
  1183 => x"5287fc80",
  1184 => x"d8519fee",
  1185 => x"2dbdac08",
  1186 => x"802e8c38",
  1187 => x"ba805185",
  1188 => x"f22d8153",
  1189 => x"a68f0481",
  1190 => x"ff0bd40c",
  1191 => x"81fe0bd4",
  1192 => x"0c80ff55",
  1193 => x"75708405",
  1194 => x"57087098",
  1195 => x"2ad40c70",
  1196 => x"902c7081",
  1197 => x"ff06d40c",
  1198 => x"5470882c",
  1199 => x"7081ff06",
  1200 => x"d40c5470",
  1201 => x"81ff06d4",
  1202 => x"0c54ff15",
  1203 => x"55748025",
  1204 => x"d33881ff",
  1205 => x"0bd40c81",
  1206 => x"ff0bd40c",
  1207 => x"81ff0bd4",
  1208 => x"0c868da0",
  1209 => x"5481ff0b",
  1210 => x"d40cd408",
  1211 => x"81ff0655",
  1212 => x"748738ff",
  1213 => x"145473ed",
  1214 => x"3881ff0b",
  1215 => x"d40cd008",
  1216 => x"708f2a70",
  1217 => x"81065151",
  1218 => x"5372f338",
  1219 => x"72d00c72",
  1220 => x"bdac0c02",
  1221 => x"98050d04",
  1222 => x"02e8050d",
  1223 => x"78558056",
  1224 => x"81ff0bd4",
  1225 => x"0cd00870",
  1226 => x"8f2a7081",
  1227 => x"06515153",
  1228 => x"72f33882",
  1229 => x"810bd00c",
  1230 => x"81ff0bd4",
  1231 => x"0c775287",
  1232 => x"fc80d151",
  1233 => x"9fee2d80",
  1234 => x"dbc6df54",
  1235 => x"bdac0880",
  1236 => x"2e8a38ba",
  1237 => x"905185f2",
  1238 => x"2da7af04",
  1239 => x"81ff0bd4",
  1240 => x"0cd40870",
  1241 => x"81ff0651",
  1242 => x"537281fe",
  1243 => x"2e098106",
  1244 => x"9d3880ff",
  1245 => x"539fa02d",
  1246 => x"bdac0875",
  1247 => x"70840557",
  1248 => x"0cff1353",
  1249 => x"728025ed",
  1250 => x"388156a7",
  1251 => x"9404ff14",
  1252 => x"5473c938",
  1253 => x"81ff0bd4",
  1254 => x"0c81ff0b",
  1255 => x"d40cd008",
  1256 => x"708f2a70",
  1257 => x"81065151",
  1258 => x"5372f338",
  1259 => x"72d00c75",
  1260 => x"bdac0c02",
  1261 => x"98050d04",
  1262 => x"02f4050d",
  1263 => x"7470882a",
  1264 => x"83fe8006",
  1265 => x"7072982a",
  1266 => x"0772882b",
  1267 => x"87fc8080",
  1268 => x"0673982b",
  1269 => x"81f00a06",
  1270 => x"71730707",
  1271 => x"bdac0c56",
  1272 => x"51535102",
  1273 => x"8c050d04",
  1274 => x"02f8050d",
  1275 => x"028e0580",
  1276 => x"f52d7488",
  1277 => x"2b077083",
  1278 => x"ffff06bd",
  1279 => x"ac0c5102",
  1280 => x"88050d04",
  1281 => x"02fc050d",
  1282 => x"72518071",
  1283 => x"0c800b84",
  1284 => x"120c0284",
  1285 => x"050d0402",
  1286 => x"f0050d75",
  1287 => x"70088412",
  1288 => x"08535353",
  1289 => x"ff547171",
  1290 => x"2ea838ab",
  1291 => x"db2d8413",
  1292 => x"08708429",
  1293 => x"14881170",
  1294 => x"087081ff",
  1295 => x"06841808",
  1296 => x"81118706",
  1297 => x"841a0c53",
  1298 => x"51555151",
  1299 => x"51abd52d",
  1300 => x"715473bd",
  1301 => x"ac0c0290",
  1302 => x"050d0402",
  1303 => x"f8050dab",
  1304 => x"db2de008",
  1305 => x"708b2a70",
  1306 => x"81065152",
  1307 => x"5270802e",
  1308 => x"a13880c7",
  1309 => x"a4087084",
  1310 => x"2980c7ac",
  1311 => x"057381ff",
  1312 => x"06710c51",
  1313 => x"5180c7a4",
  1314 => x"08811187",
  1315 => x"0680c7a4",
  1316 => x"0c51800b",
  1317 => x"80c7cc0c",
  1318 => x"abce2dab",
  1319 => x"d52d0288",
  1320 => x"050d0402",
  1321 => x"fc050dab",
  1322 => x"db2d810b",
  1323 => x"80c7cc0c",
  1324 => x"abd52d80",
  1325 => x"c7cc0851",
  1326 => x"70f93802",
  1327 => x"84050d04",
  1328 => x"02fc050d",
  1329 => x"80c7a451",
  1330 => x"a8842da8",
  1331 => x"db51abca",
  1332 => x"2daaf42d",
  1333 => x"0284050d",
  1334 => x"0402f405",
  1335 => x"0daadb04",
  1336 => x"bdac0881",
  1337 => x"f02e0981",
  1338 => x"06893881",
  1339 => x"0bbda00c",
  1340 => x"aadb04bd",
  1341 => x"ac0881e0",
  1342 => x"2e098106",
  1343 => x"8938810b",
  1344 => x"bda40caa",
  1345 => x"db04bdac",
  1346 => x"0852bda4",
  1347 => x"08802e88",
  1348 => x"38bdac08",
  1349 => x"81800552",
  1350 => x"71842c72",
  1351 => x"8f065353",
  1352 => x"bda00880",
  1353 => x"2e993872",
  1354 => x"8429bce0",
  1355 => x"05721381",
  1356 => x"712b7009",
  1357 => x"73080673",
  1358 => x"0c515353",
  1359 => x"aad10472",
  1360 => x"8429bce0",
  1361 => x"05721383",
  1362 => x"712b7208",
  1363 => x"07720c53",
  1364 => x"53800bbd",
  1365 => x"a40c800b",
  1366 => x"bda00c80",
  1367 => x"c7a451a8",
  1368 => x"972dbdac",
  1369 => x"08ff24fe",
  1370 => x"f738800b",
  1371 => x"bdac0c02",
  1372 => x"8c050d04",
  1373 => x"02f8050d",
  1374 => x"bce0528f",
  1375 => x"51807270",
  1376 => x"8405540c",
  1377 => x"ff115170",
  1378 => x"8025f238",
  1379 => x"0288050d",
  1380 => x"0402f005",
  1381 => x"0d7551ab",
  1382 => x"db2d7082",
  1383 => x"2cfc06bc",
  1384 => x"e0117210",
  1385 => x"9e067108",
  1386 => x"70722a70",
  1387 => x"83068274",
  1388 => x"2b700974",
  1389 => x"06760c54",
  1390 => x"51565753",
  1391 => x"5153abd5",
  1392 => x"2d71bdac",
  1393 => x"0c029005",
  1394 => x"0d047198",
  1395 => x"0c04ffb0",
  1396 => x"08bdac0c",
  1397 => x"04810bff",
  1398 => x"b00c0480",
  1399 => x"0bffb00c",
  1400 => x"0402fc05",
  1401 => x"0d810bbd",
  1402 => x"a80c8151",
  1403 => x"84e62d02",
  1404 => x"84050d04",
  1405 => x"02fc050d",
  1406 => x"800bbda8",
  1407 => x"0c805184",
  1408 => x"e62d0284",
  1409 => x"050d0402",
  1410 => x"ec050d76",
  1411 => x"54805287",
  1412 => x"0b881580",
  1413 => x"f52d5653",
  1414 => x"74722483",
  1415 => x"38a05372",
  1416 => x"5182ef2d",
  1417 => x"81128b15",
  1418 => x"80f52d54",
  1419 => x"52727225",
  1420 => x"de380294",
  1421 => x"050d0402",
  1422 => x"f0050d80",
  1423 => x"c7dc0854",
  1424 => x"81f82d80",
  1425 => x"0b80c7e0",
  1426 => x"0c730880",
  1427 => x"2e818438",
  1428 => x"820bbdc0",
  1429 => x"0c80c7e0",
  1430 => x"088f06bd",
  1431 => x"bc0c7308",
  1432 => x"5271832e",
  1433 => x"96387183",
  1434 => x"26893871",
  1435 => x"812eaf38",
  1436 => x"adbc0471",
  1437 => x"852e9f38",
  1438 => x"adbc0488",
  1439 => x"1480f52d",
  1440 => x"841508ba",
  1441 => x"a0535452",
  1442 => x"85f22d71",
  1443 => x"84291370",
  1444 => x"085252ad",
  1445 => x"c0047351",
  1446 => x"ac872dad",
  1447 => x"bc0480c7",
  1448 => x"d0088815",
  1449 => x"082c7081",
  1450 => x"06515271",
  1451 => x"802e8738",
  1452 => x"baa451ad",
  1453 => x"b904baa8",
  1454 => x"5185f22d",
  1455 => x"84140851",
  1456 => x"85f22d80",
  1457 => x"c7e00881",
  1458 => x"0580c7e0",
  1459 => x"0c8c1454",
  1460 => x"acc90402",
  1461 => x"90050d04",
  1462 => x"7180c7dc",
  1463 => x"0cacb72d",
  1464 => x"80c7e008",
  1465 => x"ff0580c7",
  1466 => x"e40c0402",
  1467 => x"e8050d80",
  1468 => x"c7dc0880",
  1469 => x"c7e80857",
  1470 => x"5580f851",
  1471 => x"ab912dbd",
  1472 => x"ac08812a",
  1473 => x"70810651",
  1474 => x"52719b38",
  1475 => x"8751ab91",
  1476 => x"2dbdac08",
  1477 => x"812a7081",
  1478 => x"06515271",
  1479 => x"802eb138",
  1480 => x"aea604a9",
  1481 => x"d92d8751",
  1482 => x"ab912dbd",
  1483 => x"ac08f438",
  1484 => x"aeb604a9",
  1485 => x"d92d80f8",
  1486 => x"51ab912d",
  1487 => x"bdac08f3",
  1488 => x"38bda808",
  1489 => x"813270bd",
  1490 => x"a80c7052",
  1491 => x"5284e62d",
  1492 => x"800b80c7",
  1493 => x"d40c800b",
  1494 => x"80c7d80c",
  1495 => x"bda80882",
  1496 => x"fd3880da",
  1497 => x"51ab912d",
  1498 => x"bdac0880",
  1499 => x"2e8c3880",
  1500 => x"c7d40881",
  1501 => x"800780c7",
  1502 => x"d40c80d9",
  1503 => x"51ab912d",
  1504 => x"bdac0880",
  1505 => x"2e8c3880",
  1506 => x"c7d40880",
  1507 => x"c00780c7",
  1508 => x"d40c8194",
  1509 => x"51ab912d",
  1510 => x"bdac0880",
  1511 => x"2e8b3880",
  1512 => x"c7d40890",
  1513 => x"0780c7d4",
  1514 => x"0c819151",
  1515 => x"ab912dbd",
  1516 => x"ac08802e",
  1517 => x"8b3880c7",
  1518 => x"d408a007",
  1519 => x"80c7d40c",
  1520 => x"81f551ab",
  1521 => x"912dbdac",
  1522 => x"08802e8b",
  1523 => x"3880c7d4",
  1524 => x"08810780",
  1525 => x"c7d40c81",
  1526 => x"f251ab91",
  1527 => x"2dbdac08",
  1528 => x"802e8b38",
  1529 => x"80c7d408",
  1530 => x"820780c7",
  1531 => x"d40c81eb",
  1532 => x"51ab912d",
  1533 => x"bdac0880",
  1534 => x"2e8b3880",
  1535 => x"c7d40884",
  1536 => x"0780c7d4",
  1537 => x"0c81f451",
  1538 => x"ab912dbd",
  1539 => x"ac08802e",
  1540 => x"8b3880c7",
  1541 => x"d4088807",
  1542 => x"80c7d40c",
  1543 => x"80d851ab",
  1544 => x"912dbdac",
  1545 => x"08802e8c",
  1546 => x"3880c7d8",
  1547 => x"08818007",
  1548 => x"80c7d80c",
  1549 => x"9251ab91",
  1550 => x"2dbdac08",
  1551 => x"802e8c38",
  1552 => x"80c7d808",
  1553 => x"80c00780",
  1554 => x"c7d80c94",
  1555 => x"51ab912d",
  1556 => x"bdac0880",
  1557 => x"2e8b3880",
  1558 => x"c7d80890",
  1559 => x"0780c7d8",
  1560 => x"0c9151ab",
  1561 => x"912dbdac",
  1562 => x"08802e8b",
  1563 => x"3880c7d8",
  1564 => x"08a00780",
  1565 => x"c7d80c9d",
  1566 => x"51ab912d",
  1567 => x"bdac0880",
  1568 => x"2e8b3880",
  1569 => x"c7d80881",
  1570 => x"0780c7d8",
  1571 => x"0c9b51ab",
  1572 => x"912dbdac",
  1573 => x"08802e8b",
  1574 => x"3880c7d8",
  1575 => x"08820780",
  1576 => x"c7d80c9c",
  1577 => x"51ab912d",
  1578 => x"bdac0880",
  1579 => x"2e8b3880",
  1580 => x"c7d80884",
  1581 => x"0780c7d8",
  1582 => x"0ca351ab",
  1583 => x"912dbdac",
  1584 => x"08802e8b",
  1585 => x"3880c7d8",
  1586 => x"08880780",
  1587 => x"c7d80c81",
  1588 => x"fd51ab91",
  1589 => x"2d81fa51",
  1590 => x"ab912db7",
  1591 => x"a60481f5",
  1592 => x"51ab912d",
  1593 => x"bdac0881",
  1594 => x"2a708106",
  1595 => x"51527180",
  1596 => x"2eb33880",
  1597 => x"c7e40852",
  1598 => x"71802e8a",
  1599 => x"38ff1280",
  1600 => x"c7e40cb2",
  1601 => x"a50480c7",
  1602 => x"e0081080",
  1603 => x"c7e00805",
  1604 => x"70842916",
  1605 => x"51528812",
  1606 => x"08802e89",
  1607 => x"38ff5188",
  1608 => x"12085271",
  1609 => x"2d81f251",
  1610 => x"ab912dbd",
  1611 => x"ac08812a",
  1612 => x"70810651",
  1613 => x"5271802e",
  1614 => x"b43880c7",
  1615 => x"e008ff11",
  1616 => x"80c7e408",
  1617 => x"56535373",
  1618 => x"72258a38",
  1619 => x"811480c7",
  1620 => x"e40cb2ed",
  1621 => x"04721013",
  1622 => x"70842916",
  1623 => x"51528812",
  1624 => x"08802e89",
  1625 => x"38fe5188",
  1626 => x"12085271",
  1627 => x"2d81fd51",
  1628 => x"ab912dbd",
  1629 => x"ac08812a",
  1630 => x"70810651",
  1631 => x"5271802e",
  1632 => x"b13880c7",
  1633 => x"e408802e",
  1634 => x"8a38800b",
  1635 => x"80c7e40c",
  1636 => x"b3b20480",
  1637 => x"c7e00810",
  1638 => x"80c7e008",
  1639 => x"05708429",
  1640 => x"16515288",
  1641 => x"1208802e",
  1642 => x"8938fd51",
  1643 => x"88120852",
  1644 => x"712d81fa",
  1645 => x"51ab912d",
  1646 => x"bdac0881",
  1647 => x"2a708106",
  1648 => x"51527180",
  1649 => x"2eb13880",
  1650 => x"c7e008ff",
  1651 => x"11545280",
  1652 => x"c7e40873",
  1653 => x"25893872",
  1654 => x"80c7e40c",
  1655 => x"b3f70471",
  1656 => x"10127084",
  1657 => x"29165152",
  1658 => x"88120880",
  1659 => x"2e8938fc",
  1660 => x"51881208",
  1661 => x"52712d80",
  1662 => x"c7e40870",
  1663 => x"53547380",
  1664 => x"2e8a388c",
  1665 => x"15ff1555",
  1666 => x"55b3fe04",
  1667 => x"820bbdc0",
  1668 => x"0c718f06",
  1669 => x"bdbc0c81",
  1670 => x"eb51ab91",
  1671 => x"2dbdac08",
  1672 => x"812a7081",
  1673 => x"06515271",
  1674 => x"802ead38",
  1675 => x"7408852e",
  1676 => x"098106a4",
  1677 => x"38881580",
  1678 => x"f52dff05",
  1679 => x"52718816",
  1680 => x"81b72d71",
  1681 => x"982b5271",
  1682 => x"80258838",
  1683 => x"800b8816",
  1684 => x"81b72d74",
  1685 => x"51ac872d",
  1686 => x"81f451ab",
  1687 => x"912dbdac",
  1688 => x"08812a70",
  1689 => x"81065152",
  1690 => x"71802eb3",
  1691 => x"38740885",
  1692 => x"2e098106",
  1693 => x"aa388815",
  1694 => x"80f52d81",
  1695 => x"05527188",
  1696 => x"1681b72d",
  1697 => x"7181ff06",
  1698 => x"8b1680f5",
  1699 => x"2d545272",
  1700 => x"72278738",
  1701 => x"72881681",
  1702 => x"b72d7451",
  1703 => x"ac872d80",
  1704 => x"da51ab91",
  1705 => x"2dbdac08",
  1706 => x"812a7081",
  1707 => x"06515271",
  1708 => x"802e81ac",
  1709 => x"3880c7dc",
  1710 => x"0880c7e4",
  1711 => x"08555373",
  1712 => x"802e8a38",
  1713 => x"8c13ff15",
  1714 => x"5553b5bf",
  1715 => x"04720852",
  1716 => x"71822ea6",
  1717 => x"38718226",
  1718 => x"89387181",
  1719 => x"2eaa38b6",
  1720 => x"e0047183",
  1721 => x"2eb43871",
  1722 => x"842e0981",
  1723 => x"0680f138",
  1724 => x"88130851",
  1725 => x"add82db6",
  1726 => x"e00480c7",
  1727 => x"e4085188",
  1728 => x"13085271",
  1729 => x"2db6e004",
  1730 => x"810b8814",
  1731 => x"082b80c7",
  1732 => x"d0083280",
  1733 => x"c7d00cb6",
  1734 => x"b5048813",
  1735 => x"80f52d81",
  1736 => x"058b1480",
  1737 => x"f52d5354",
  1738 => x"71742483",
  1739 => x"38805473",
  1740 => x"881481b7",
  1741 => x"2dacb72d",
  1742 => x"b6e00475",
  1743 => x"08802ea3",
  1744 => x"38750851",
  1745 => x"ab912dbd",
  1746 => x"ac088106",
  1747 => x"5271802e",
  1748 => x"8c3880c7",
  1749 => x"e4085184",
  1750 => x"16085271",
  1751 => x"2d881656",
  1752 => x"75d93880",
  1753 => x"54800bbd",
  1754 => x"c00c738f",
  1755 => x"06bdbc0c",
  1756 => x"a0527380",
  1757 => x"c7e4082e",
  1758 => x"09810699",
  1759 => x"3880c7e0",
  1760 => x"08ff0574",
  1761 => x"32700981",
  1762 => x"05707207",
  1763 => x"9f2a9171",
  1764 => x"31515153",
  1765 => x"53715182",
  1766 => x"ef2d8114",
  1767 => x"548e7425",
  1768 => x"c438bda8",
  1769 => x"085271bd",
  1770 => x"ac0c0298",
  1771 => x"050d0400",
  1772 => x"00ffffff",
  1773 => x"ff00ffff",
  1774 => x"ffff00ff",
  1775 => x"ffffff00",
  1776 => x"52657365",
  1777 => x"74000000",
  1778 => x"53617665",
  1779 => x"20736574",
  1780 => x"74696e67",
  1781 => x"73000000",
  1782 => x"5363616e",
  1783 => x"6c696e65",
  1784 => x"73000000",
  1785 => x"4c6f6164",
  1786 => x"20524f4d",
  1787 => x"20100000",
  1788 => x"45786974",
  1789 => x"00000000",
  1790 => x"4a6f7973",
  1791 => x"7469636b",
  1792 => x"20737761",
  1793 => x"70000000",
  1794 => x"4a6f7973",
  1795 => x"7469636b",
  1796 => x"206e6f72",
  1797 => x"6d616c00",
  1798 => x"56474120",
  1799 => x"2d203331",
  1800 => x"4b487a2c",
  1801 => x"20363048",
  1802 => x"7a000000",
  1803 => x"5456202d",
  1804 => x"20343830",
  1805 => x"692c2036",
  1806 => x"30487a00",
  1807 => x"4261636b",
  1808 => x"00000000",
  1809 => x"46504741",
  1810 => x"47454e20",
  1811 => x"43464700",
  1812 => x"496e6974",
  1813 => x"69616c69",
  1814 => x"7a696e67",
  1815 => x"20534420",
  1816 => x"63617264",
  1817 => x"0a000000",
  1818 => x"424f4f54",
  1819 => x"20202020",
  1820 => x"47454e00",
  1821 => x"43617264",
  1822 => x"20696e69",
  1823 => x"74206661",
  1824 => x"696c6564",
  1825 => x"0a000000",
  1826 => x"4d425220",
  1827 => x"6661696c",
  1828 => x"0a000000",
  1829 => x"46415431",
  1830 => x"36202020",
  1831 => x"00000000",
  1832 => x"46415433",
  1833 => x"32202020",
  1834 => x"00000000",
  1835 => x"4e6f2070",
  1836 => x"61727469",
  1837 => x"74696f6e",
  1838 => x"20736967",
  1839 => x"0a000000",
  1840 => x"42616420",
  1841 => x"70617274",
  1842 => x"0a000000",
  1843 => x"53444843",
  1844 => x"20657272",
  1845 => x"6f72210a",
  1846 => x"00000000",
  1847 => x"53442069",
  1848 => x"6e69742e",
  1849 => x"2e2e0a00",
  1850 => x"53442063",
  1851 => x"61726420",
  1852 => x"72657365",
  1853 => x"74206661",
  1854 => x"696c6564",
  1855 => x"210a0000",
  1856 => x"57726974",
  1857 => x"65206661",
  1858 => x"696c6564",
  1859 => x"0a000000",
  1860 => x"52656164",
  1861 => x"20666169",
  1862 => x"6c65640a",
  1863 => x"00000000",
  1864 => x"16200000",
  1865 => x"14200000",
  1866 => x"15200000",
  1867 => x"00000002",
  1868 => x"00000000",
  1869 => x"00000002",
  1870 => x"00001bc0",
  1871 => x"000004aa",
  1872 => x"00000002",
  1873 => x"00001bc8",
  1874 => x"0000037d",
  1875 => x"00000003",
  1876 => x"00001d9c",
  1877 => x"00000002",
  1878 => x"00000001",
  1879 => x"00001bd8",
  1880 => x"00000001",
  1881 => x"00000003",
  1882 => x"00001d94",
  1883 => x"00000002",
  1884 => x"00000002",
  1885 => x"00001be4",
  1886 => x"00000744",
  1887 => x"00000002",
  1888 => x"00001bf0",
  1889 => x"000015f4",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00001bf8",
  1894 => x"00001c08",
  1895 => x"00001c18",
  1896 => x"00001c2c",
  1897 => x"00000002",
  1898 => x"00001edc",
  1899 => x"00000538",
  1900 => x"00000002",
  1901 => x"00001efa",
  1902 => x"00000538",
  1903 => x"00000002",
  1904 => x"00001f18",
  1905 => x"00000538",
  1906 => x"00000002",
  1907 => x"00001f36",
  1908 => x"00000538",
  1909 => x"00000002",
  1910 => x"00001f54",
  1911 => x"00000538",
  1912 => x"00000002",
  1913 => x"00001f72",
  1914 => x"00000538",
  1915 => x"00000002",
  1916 => x"00001f90",
  1917 => x"00000538",
  1918 => x"00000002",
  1919 => x"00001fae",
  1920 => x"00000538",
  1921 => x"00000002",
  1922 => x"00001fcc",
  1923 => x"00000538",
  1924 => x"00000002",
  1925 => x"00001fea",
  1926 => x"00000538",
  1927 => x"00000002",
  1928 => x"00002008",
  1929 => x"00000538",
  1930 => x"00000002",
  1931 => x"00002026",
  1932 => x"00000538",
  1933 => x"00000002",
  1934 => x"00002044",
  1935 => x"00000538",
  1936 => x"00000004",
  1937 => x"00001c3c",
  1938 => x"00001d34",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"000006d8",
  1942 => x"00000000",
  1943 => x"00000000",
  1944 => x"00000000",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

