-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbc",
     9 => x"d8080b0b",
    10 => x"0bbcdc08",
    11 => x"0b0b0bbc",
    12 => x"e0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bce00c0b",
    16 => x"0b0bbcdc",
    17 => x"0c0b0b0b",
    18 => x"bcd80c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb790",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bcd87080",
    57 => x"c798278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518efa04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbce80c",
    65 => x"9f0bbcec",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bcec08ff",
    69 => x"05bcec0c",
    70 => x"bcec0880",
    71 => x"25eb38bc",
    72 => x"e808ff05",
    73 => x"bce80cbc",
    74 => x"e8088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbc",
    94 => x"e808258f",
    95 => x"3882b32d",
    96 => x"bce808ff",
    97 => x"05bce80c",
    98 => x"82f504bc",
    99 => x"e808bcec",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038bce8",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"bcec0881",
   109 => x"05bcec0c",
   110 => x"bcec0851",
   111 => x"9f7125e2",
   112 => x"38800bbc",
   113 => x"ec0cbce8",
   114 => x"088105bc",
   115 => x"e80c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34bcec08",
   120 => x"8105bcec",
   121 => x"0cbcec08",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbcec0c",
   125 => x"bce80881",
   126 => x"05bce80c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"bcf00cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbc",
   162 => x"f00c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72bcf008",
   167 => x"8407bcf0",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"b9ec0c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"bcf00852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"fc050d72",
   198 => x"70820680",
   199 => x"c6fc0c70",
   200 => x"81065151",
   201 => x"70ba940b",
   202 => x"81b72d70",
   203 => x"bcd80c02",
   204 => x"84050d04",
   205 => x"02f8050d",
   206 => x"b88452bc",
   207 => x"f4519bed",
   208 => x"2dbcd808",
   209 => x"802ea138",
   210 => x"80c09052",
   211 => x"bcf4519e",
   212 => x"ae2d80c0",
   213 => x"9008bd80",
   214 => x"0c80c090",
   215 => x"08fec00c",
   216 => x"80c09008",
   217 => x"5186932d",
   218 => x"0288050d",
   219 => x"0402f005",
   220 => x"0d805191",
   221 => x"bc2db884",
   222 => x"52bcf451",
   223 => x"9bed2dbc",
   224 => x"d808802e",
   225 => x"a838bd80",
   226 => x"0880c090",
   227 => x"0c80c094",
   228 => x"5480fd53",
   229 => x"80747084",
   230 => x"05560cff",
   231 => x"13537280",
   232 => x"25f23880",
   233 => x"c09052bc",
   234 => x"f4519ed7",
   235 => x"2d029005",
   236 => x"0d0402d8",
   237 => x"050d800b",
   238 => x"b9f00cbd",
   239 => x"8008fec0",
   240 => x"0c810bfe",
   241 => x"c40c840b",
   242 => x"fec40c7b",
   243 => x"52bcf451",
   244 => x"9bed2dbc",
   245 => x"d80853bc",
   246 => x"d808802e",
   247 => x"81b338bc",
   248 => x"f8085580",
   249 => x"0bff1657",
   250 => x"5975792e",
   251 => x"8b388119",
   252 => x"76812a57",
   253 => x"5975f738",
   254 => x"f7195974",
   255 => x"b080802e",
   256 => x"09810689",
   257 => x"38820bfe",
   258 => x"dc0c88a4",
   259 => x"04749880",
   260 => x"802e0981",
   261 => x"06893881",
   262 => x"0bfedc0c",
   263 => x"88a40480",
   264 => x"0bfedc0c",
   265 => x"815a8075",
   266 => x"2580df38",
   267 => x"78527551",
   268 => x"84812d80",
   269 => x"c09052bc",
   270 => x"f4519eae",
   271 => x"2dbcd808",
   272 => x"802ea838",
   273 => x"80c09058",
   274 => x"83fc5777",
   275 => x"70840559",
   276 => x"087083ff",
   277 => x"ff067190",
   278 => x"2afec80c",
   279 => x"fec80cfc",
   280 => x"18585376",
   281 => x"8025e438",
   282 => x"88f204bc",
   283 => x"d8085a84",
   284 => x"8055bcf4",
   285 => x"519e802d",
   286 => x"fc801581",
   287 => x"17575574",
   288 => x"8024ffa8",
   289 => x"3879802e",
   290 => x"8638820b",
   291 => x"b9f00c79",
   292 => x"5372bcd8",
   293 => x"0c02a805",
   294 => x"0d0402fc",
   295 => x"050dabd4",
   296 => x"2dfec451",
   297 => x"81710c82",
   298 => x"710c0284",
   299 => x"050d0402",
   300 => x"f4050d74",
   301 => x"76785354",
   302 => x"52807125",
   303 => x"97387270",
   304 => x"81055480",
   305 => x"f52d7270",
   306 => x"81055481",
   307 => x"b72dff11",
   308 => x"5170eb38",
   309 => x"807281b7",
   310 => x"2d028c05",
   311 => x"0d0402e8",
   312 => x"050d7756",
   313 => x"80705654",
   314 => x"737624b3",
   315 => x"3880c6a0",
   316 => x"08742eab",
   317 => x"38735199",
   318 => x"b62dbcd8",
   319 => x"08bcd808",
   320 => x"09810570",
   321 => x"bcd80807",
   322 => x"9f2a7705",
   323 => x"81175757",
   324 => x"53537476",
   325 => x"24893880",
   326 => x"c6a00874",
   327 => x"26d73872",
   328 => x"bcd80c02",
   329 => x"98050d04",
   330 => x"02f4050d",
   331 => x"bc840815",
   332 => x"5189de2d",
   333 => x"bcd80880",
   334 => x"2e95388b",
   335 => x"53bcd808",
   336 => x"5280c490",
   337 => x"5189af2d",
   338 => x"80c49051",
   339 => x"87b22db9",
   340 => x"f451adb8",
   341 => x"2dabd42d",
   342 => x"805184e6",
   343 => x"2d028c05",
   344 => x"0d0402dc",
   345 => x"050d8070",
   346 => x"5a5574bc",
   347 => x"840825b1",
   348 => x"3880c6a0",
   349 => x"08752ea9",
   350 => x"38785199",
   351 => x"b62dbcd8",
   352 => x"08098105",
   353 => x"70bcd808",
   354 => x"079f2a76",
   355 => x"05811b5b",
   356 => x"565474bc",
   357 => x"84082589",
   358 => x"3880c6a0",
   359 => x"087926d9",
   360 => x"38805578",
   361 => x"80c6a008",
   362 => x"2781d038",
   363 => x"785199b6",
   364 => x"2dbcd808",
   365 => x"802e81a5",
   366 => x"38bcd808",
   367 => x"8b0580f5",
   368 => x"2d70842a",
   369 => x"70810677",
   370 => x"1078842b",
   371 => x"80c4900b",
   372 => x"80f52d5c",
   373 => x"5c535155",
   374 => x"5673802e",
   375 => x"80c73874",
   376 => x"16822b8d",
   377 => x"9e0bbad8",
   378 => x"120c5477",
   379 => x"753110bd",
   380 => x"88115556",
   381 => x"90747081",
   382 => x"055681b7",
   383 => x"2da07481",
   384 => x"b72d7681",
   385 => x"ff068116",
   386 => x"58547380",
   387 => x"2e8a389c",
   388 => x"5380c490",
   389 => x"528c9e04",
   390 => x"8b53bcd8",
   391 => x"0852bd8a",
   392 => x"16518cd5",
   393 => x"04741682",
   394 => x"2b8aa80b",
   395 => x"bad8120c",
   396 => x"547681ff",
   397 => x"06811658",
   398 => x"5473802e",
   399 => x"8a389c53",
   400 => x"80c49052",
   401 => x"8ccd048b",
   402 => x"53bcd808",
   403 => x"52777531",
   404 => x"10bd8805",
   405 => x"51765589",
   406 => x"af2d8cf0",
   407 => x"04749029",
   408 => x"75317010",
   409 => x"bd880551",
   410 => x"54bcd808",
   411 => x"7481b72d",
   412 => x"81195974",
   413 => x"8b24a238",
   414 => x"8ba30474",
   415 => x"90297531",
   416 => x"7010bd88",
   417 => x"058c7731",
   418 => x"57515480",
   419 => x"7481b72d",
   420 => x"9e14ff16",
   421 => x"565474f3",
   422 => x"3802a405",
   423 => x"0d0402fc",
   424 => x"050dbc84",
   425 => x"08135189",
   426 => x"de2dbcd8",
   427 => x"08802e88",
   428 => x"38bcd808",
   429 => x"5191bc2d",
   430 => x"800bbc84",
   431 => x"0c8ae22d",
   432 => x"ac972d02",
   433 => x"84050d04",
   434 => x"02fc050d",
   435 => x"725170fd",
   436 => x"2ead3870",
   437 => x"fd248a38",
   438 => x"70fc2e80",
   439 => x"c4388ea9",
   440 => x"0470fe2e",
   441 => x"b13870ff",
   442 => x"2e098106",
   443 => x"bc38bc84",
   444 => x"08517080",
   445 => x"2eb338ff",
   446 => x"11bc840c",
   447 => x"8ea904bc",
   448 => x"8408f005",
   449 => x"70bc840c",
   450 => x"51708025",
   451 => x"9c38800b",
   452 => x"bc840c8e",
   453 => x"a904bc84",
   454 => x"088105bc",
   455 => x"840c8ea9",
   456 => x"04bc8408",
   457 => x"9005bc84",
   458 => x"0c8ae22d",
   459 => x"ac972d02",
   460 => x"84050d04",
   461 => x"02fc050d",
   462 => x"800bbc84",
   463 => x"0c8ae22d",
   464 => x"bad051ad",
   465 => x"b82d0284",
   466 => x"050d0402",
   467 => x"f8050d80",
   468 => x"c6fc0882",
   469 => x"06ba940b",
   470 => x"80f52d52",
   471 => x"5270802e",
   472 => x"85387181",
   473 => x"0752bd84",
   474 => x"08802e85",
   475 => x"38719007",
   476 => x"5271bcd8",
   477 => x"0c028805",
   478 => x"0d0402f4",
   479 => x"050d810b",
   480 => x"bd840c80",
   481 => x"0bb9f00c",
   482 => x"90518693",
   483 => x"2d810bfe",
   484 => x"c40c840b",
   485 => x"fec40c83",
   486 => x"0bfecc0c",
   487 => x"b8905185",
   488 => x"f22d8452",
   489 => x"a38e2d92",
   490 => x"dd2dbcd8",
   491 => x"08802e86",
   492 => x"38fe528f",
   493 => x"be04ff12",
   494 => x"52718024",
   495 => x"e7387180",
   496 => x"2e81ab38",
   497 => x"a9a02dab",
   498 => x"b52da983",
   499 => x"2da9832d",
   500 => x"81f82d81",
   501 => x"5184e62d",
   502 => x"a9832da9",
   503 => x"832d8151",
   504 => x"84e62d86",
   505 => x"b42db8a8",
   506 => x"5187b22d",
   507 => x"bcd80880",
   508 => x"2e9438b9",
   509 => x"f451adb8",
   510 => x"2d805184",
   511 => x"e62d820b",
   512 => x"b9f00c90",
   513 => x"9004bcd8",
   514 => x"08518eb4",
   515 => x"2dabc12d",
   516 => x"a9b92dad",
   517 => x"cb2dbcd8",
   518 => x"0880c780",
   519 => x"08882b80",
   520 => x"c7840807",
   521 => x"fed80c53",
   522 => x"8ecb2dbc",
   523 => x"d808bd80",
   524 => x"082ea238",
   525 => x"bcd808bd",
   526 => x"800cbcd8",
   527 => x"08fec00c",
   528 => x"84527251",
   529 => x"84e62da9",
   530 => x"832da983",
   531 => x"2dff1252",
   532 => x"718025ee",
   533 => x"3872802e",
   534 => x"8c38b9f0",
   535 => x"088807fe",
   536 => x"c40c9090",
   537 => x"04b9f008",
   538 => x"fec40c90",
   539 => x"9004b8b4",
   540 => x"5185f22d",
   541 => x"800bbcd8",
   542 => x"0c028c05",
   543 => x"0d0402e8",
   544 => x"050d7779",
   545 => x"7b585555",
   546 => x"80537276",
   547 => x"25a33874",
   548 => x"70810556",
   549 => x"80f52d74",
   550 => x"70810556",
   551 => x"80f52d52",
   552 => x"5271712e",
   553 => x"86388151",
   554 => x"91b30481",
   555 => x"1353918a",
   556 => x"04805170",
   557 => x"bcd80c02",
   558 => x"98050d04",
   559 => x"02ec050d",
   560 => x"76557480",
   561 => x"2ebe389a",
   562 => x"1580e02d",
   563 => x"51a7c82d",
   564 => x"bcd808bc",
   565 => x"d80880c6",
   566 => x"c00cbcd8",
   567 => x"08545480",
   568 => x"c69c0880",
   569 => x"2e993894",
   570 => x"1580e02d",
   571 => x"51a7c82d",
   572 => x"bcd80890",
   573 => x"2b83fff0",
   574 => x"0a067075",
   575 => x"07515372",
   576 => x"80c6c00c",
   577 => x"80c6c008",
   578 => x"5372802e",
   579 => x"9d3880c6",
   580 => x"9408fe14",
   581 => x"712980c6",
   582 => x"a8080580",
   583 => x"c6c40c70",
   584 => x"842b80c6",
   585 => x"a00c5492",
   586 => x"d80480c6",
   587 => x"ac0880c6",
   588 => x"c00c80c6",
   589 => x"b00880c6",
   590 => x"c40c80c6",
   591 => x"9c08802e",
   592 => x"8b3880c6",
   593 => x"9408842b",
   594 => x"5392d304",
   595 => x"80c6b408",
   596 => x"842b5372",
   597 => x"80c6a00c",
   598 => x"0294050d",
   599 => x"0402d805",
   600 => x"0d800b80",
   601 => x"c69c0c80",
   602 => x"c0905280",
   603 => x"51a5f82d",
   604 => x"bcd80854",
   605 => x"bcd8088c",
   606 => x"38b8c851",
   607 => x"85f22d73",
   608 => x"5598b904",
   609 => x"8056810b",
   610 => x"80c6c80c",
   611 => x"8853b8d4",
   612 => x"5280c0c6",
   613 => x"5190fe2d",
   614 => x"bcd80876",
   615 => x"2e098106",
   616 => x"8838bcd8",
   617 => x"0880c6c8",
   618 => x"0c8853b8",
   619 => x"e05280c0",
   620 => x"e25190fe",
   621 => x"2dbcd808",
   622 => x"8838bcd8",
   623 => x"0880c6c8",
   624 => x"0c80c6c8",
   625 => x"08802e80",
   626 => x"fd3880c3",
   627 => x"d60b80f5",
   628 => x"2d80c3d7",
   629 => x"0b80f52d",
   630 => x"71982b71",
   631 => x"902b0780",
   632 => x"c3d80b80",
   633 => x"f52d7088",
   634 => x"2b720780",
   635 => x"c3d90b80",
   636 => x"f52d7107",
   637 => x"80c48e0b",
   638 => x"80f52d80",
   639 => x"c48f0b80",
   640 => x"f52d7188",
   641 => x"2b07535f",
   642 => x"54525a56",
   643 => x"57557381",
   644 => x"abaa2e09",
   645 => x"81068d38",
   646 => x"7551a798",
   647 => x"2dbcd808",
   648 => x"5694b104",
   649 => x"7382d4d5",
   650 => x"2e8738b8",
   651 => x"ec5194f6",
   652 => x"0480c090",
   653 => x"527551a5",
   654 => x"f82dbcd8",
   655 => x"0855bcd8",
   656 => x"08802e83",
   657 => x"f4388853",
   658 => x"b8e05280",
   659 => x"c0e25190",
   660 => x"fe2dbcd8",
   661 => x"088a3881",
   662 => x"0b80c69c",
   663 => x"0c94fc04",
   664 => x"8853b8d4",
   665 => x"5280c0c6",
   666 => x"5190fe2d",
   667 => x"bcd80880",
   668 => x"2e8a38b9",
   669 => x"805185f2",
   670 => x"2d95db04",
   671 => x"80c48e0b",
   672 => x"80f52d54",
   673 => x"7380d52e",
   674 => x"09810680",
   675 => x"ce3880c4",
   676 => x"8f0b80f5",
   677 => x"2d547381",
   678 => x"aa2e0981",
   679 => x"06bd3880",
   680 => x"0b80c090",
   681 => x"0b80f52d",
   682 => x"56547481",
   683 => x"e92e8338",
   684 => x"81547481",
   685 => x"eb2e8c38",
   686 => x"80557375",
   687 => x"2e098106",
   688 => x"82f73880",
   689 => x"c09b0b80",
   690 => x"f52d5574",
   691 => x"8e3880c0",
   692 => x"9c0b80f5",
   693 => x"2d547382",
   694 => x"2e863880",
   695 => x"5598b904",
   696 => x"80c09d0b",
   697 => x"80f52d70",
   698 => x"80c6940c",
   699 => x"ff0580c6",
   700 => x"980c80c0",
   701 => x"9e0b80f5",
   702 => x"2d80c09f",
   703 => x"0b80f52d",
   704 => x"58760577",
   705 => x"82802905",
   706 => x"7080c6a4",
   707 => x"0c80c0a0",
   708 => x"0b80f52d",
   709 => x"7080c6b8",
   710 => x"0c80c69c",
   711 => x"08595758",
   712 => x"76802e81",
   713 => x"b5388853",
   714 => x"b8e05280",
   715 => x"c0e25190",
   716 => x"fe2dbcd8",
   717 => x"08828238",
   718 => x"80c69408",
   719 => x"70842b80",
   720 => x"c6a00c70",
   721 => x"80c6b40c",
   722 => x"80c0b50b",
   723 => x"80f52d80",
   724 => x"c0b40b80",
   725 => x"f52d7182",
   726 => x"80290580",
   727 => x"c0b60b80",
   728 => x"f52d7084",
   729 => x"80802912",
   730 => x"80c0b70b",
   731 => x"80f52d70",
   732 => x"81800a29",
   733 => x"127080c6",
   734 => x"bc0c80c6",
   735 => x"b8087129",
   736 => x"80c6a408",
   737 => x"057080c6",
   738 => x"a80c80c0",
   739 => x"bd0b80f5",
   740 => x"2d80c0bc",
   741 => x"0b80f52d",
   742 => x"71828029",
   743 => x"0580c0be",
   744 => x"0b80f52d",
   745 => x"70848080",
   746 => x"291280c0",
   747 => x"bf0b80f5",
   748 => x"2d70982b",
   749 => x"81f00a06",
   750 => x"72057080",
   751 => x"c6ac0cfe",
   752 => x"117e2977",
   753 => x"0580c6b0",
   754 => x"0c525952",
   755 => x"43545e51",
   756 => x"5259525d",
   757 => x"57595798",
   758 => x"b20480c0",
   759 => x"a20b80f5",
   760 => x"2d80c0a1",
   761 => x"0b80f52d",
   762 => x"71828029",
   763 => x"057080c6",
   764 => x"a00c70a0",
   765 => x"2983ff05",
   766 => x"70892a70",
   767 => x"80c6b40c",
   768 => x"80c0a70b",
   769 => x"80f52d80",
   770 => x"c0a60b80",
   771 => x"f52d7182",
   772 => x"80290570",
   773 => x"80c6bc0c",
   774 => x"7b71291e",
   775 => x"7080c6b0",
   776 => x"0c7d80c6",
   777 => x"ac0c7305",
   778 => x"80c6a80c",
   779 => x"555e5151",
   780 => x"55558051",
   781 => x"91bc2d81",
   782 => x"5574bcd8",
   783 => x"0c02a805",
   784 => x"0d0402ec",
   785 => x"050d7670",
   786 => x"872c7180",
   787 => x"ff065556",
   788 => x"5480c69c",
   789 => x"088a3873",
   790 => x"882c7481",
   791 => x"ff065455",
   792 => x"80c09052",
   793 => x"80c6a408",
   794 => x"1551a5f8",
   795 => x"2dbcd808",
   796 => x"54bcd808",
   797 => x"802eb638",
   798 => x"80c69c08",
   799 => x"802e9938",
   800 => x"72842980",
   801 => x"c0900570",
   802 => x"085253a7",
   803 => x"982dbcd8",
   804 => x"08f00a06",
   805 => x"5399ab04",
   806 => x"721080c0",
   807 => x"90057080",
   808 => x"e02d5253",
   809 => x"a7c82dbc",
   810 => x"d8085372",
   811 => x"5473bcd8",
   812 => x"0c029405",
   813 => x"0d0402e0",
   814 => x"050d7970",
   815 => x"842c80c6",
   816 => x"c4080571",
   817 => x"8f065255",
   818 => x"53728a38",
   819 => x"80c09052",
   820 => x"7351a5f8",
   821 => x"2d72a029",
   822 => x"80c09005",
   823 => x"54807480",
   824 => x"f52d5653",
   825 => x"74732e83",
   826 => x"38815374",
   827 => x"81e52e81",
   828 => x"f1388170",
   829 => x"74065458",
   830 => x"72802e81",
   831 => x"e5388b14",
   832 => x"80f52d70",
   833 => x"832a7906",
   834 => x"58567699",
   835 => x"38bc8808",
   836 => x"53728938",
   837 => x"7280c490",
   838 => x"0b81b72d",
   839 => x"76bc880c",
   840 => x"73539be4",
   841 => x"04758f2e",
   842 => x"09810681",
   843 => x"b538749f",
   844 => x"068d2980",
   845 => x"c4831151",
   846 => x"53811480",
   847 => x"f52d7370",
   848 => x"81055581",
   849 => x"b72d8314",
   850 => x"80f52d73",
   851 => x"70810555",
   852 => x"81b72d85",
   853 => x"1480f52d",
   854 => x"73708105",
   855 => x"5581b72d",
   856 => x"871480f5",
   857 => x"2d737081",
   858 => x"055581b7",
   859 => x"2d891480",
   860 => x"f52d7370",
   861 => x"81055581",
   862 => x"b72d8e14",
   863 => x"80f52d73",
   864 => x"70810555",
   865 => x"81b72d90",
   866 => x"1480f52d",
   867 => x"73708105",
   868 => x"5581b72d",
   869 => x"921480f5",
   870 => x"2d737081",
   871 => x"055581b7",
   872 => x"2d941480",
   873 => x"f52d7370",
   874 => x"81055581",
   875 => x"b72d9614",
   876 => x"80f52d73",
   877 => x"70810555",
   878 => x"81b72d98",
   879 => x"1480f52d",
   880 => x"73708105",
   881 => x"5581b72d",
   882 => x"9c1480f5",
   883 => x"2d737081",
   884 => x"055581b7",
   885 => x"2d9e1480",
   886 => x"f52d7381",
   887 => x"b72d77bc",
   888 => x"880c8053",
   889 => x"72bcd80c",
   890 => x"02a0050d",
   891 => x"0402cc05",
   892 => x"0d7e605e",
   893 => x"5a800b80",
   894 => x"c6c00880",
   895 => x"c6c40859",
   896 => x"5c568058",
   897 => x"80c6a008",
   898 => x"782e81b2",
   899 => x"38778f06",
   900 => x"a0175754",
   901 => x"73913880",
   902 => x"c0905276",
   903 => x"51811757",
   904 => x"a5f82d80",
   905 => x"c0905680",
   906 => x"7680f52d",
   907 => x"56547474",
   908 => x"2e833881",
   909 => x"547481e5",
   910 => x"2e80f738",
   911 => x"81707506",
   912 => x"555c7380",
   913 => x"2e80eb38",
   914 => x"8b1680f5",
   915 => x"2d980659",
   916 => x"7880df38",
   917 => x"8b537c52",
   918 => x"755190fe",
   919 => x"2dbcd808",
   920 => x"80d0389c",
   921 => x"160851a7",
   922 => x"982dbcd8",
   923 => x"08841b0c",
   924 => x"9a1680e0",
   925 => x"2d51a7c8",
   926 => x"2dbcd808",
   927 => x"bcd80888",
   928 => x"1c0cbcd8",
   929 => x"08555580",
   930 => x"c69c0880",
   931 => x"2e983894",
   932 => x"1680e02d",
   933 => x"51a7c82d",
   934 => x"bcd80890",
   935 => x"2b83fff0",
   936 => x"0a067016",
   937 => x"51547388",
   938 => x"1b0c787a",
   939 => x"0c7b549d",
   940 => x"f7048118",
   941 => x"5880c6a0",
   942 => x"087826fe",
   943 => x"d03880c6",
   944 => x"9c08802e",
   945 => x"b0387a51",
   946 => x"98c22dbc",
   947 => x"d808bcd8",
   948 => x"0880ffff",
   949 => x"fff80655",
   950 => x"5b7380ff",
   951 => x"fffff82e",
   952 => x"9438bcd8",
   953 => x"08fe0580",
   954 => x"c6940829",
   955 => x"80c6a808",
   956 => x"05579c82",
   957 => x"04805473",
   958 => x"bcd80c02",
   959 => x"b4050d04",
   960 => x"02f4050d",
   961 => x"74700881",
   962 => x"05710c70",
   963 => x"0880c698",
   964 => x"08065353",
   965 => x"718e3888",
   966 => x"13085198",
   967 => x"c22dbcd8",
   968 => x"0888140c",
   969 => x"810bbcd8",
   970 => x"0c028c05",
   971 => x"0d0402f0",
   972 => x"050d7588",
   973 => x"1108fe05",
   974 => x"80c69408",
   975 => x"2980c6a8",
   976 => x"08117208",
   977 => x"80c69808",
   978 => x"06057955",
   979 => x"535454a5",
   980 => x"f82d0290",
   981 => x"050d0402",
   982 => x"f0050d75",
   983 => x"881108fe",
   984 => x"0580c694",
   985 => x"082980c6",
   986 => x"a8081172",
   987 => x"0880c698",
   988 => x"08060579",
   989 => x"55535454",
   990 => x"a4b82d02",
   991 => x"90050d04",
   992 => x"02f4050d",
   993 => x"d45281ff",
   994 => x"720c7108",
   995 => x"5381ff72",
   996 => x"0c72882b",
   997 => x"83fe8006",
   998 => x"72087081",
   999 => x"ff065152",
  1000 => x"5381ff72",
  1001 => x"0c727107",
  1002 => x"882b7208",
  1003 => x"7081ff06",
  1004 => x"51525381",
  1005 => x"ff720c72",
  1006 => x"7107882b",
  1007 => x"72087081",
  1008 => x"ff067207",
  1009 => x"bcd80c52",
  1010 => x"53028c05",
  1011 => x"0d0402f4",
  1012 => x"050d7476",
  1013 => x"7181ff06",
  1014 => x"d40c5353",
  1015 => x"80c6cc08",
  1016 => x"85387189",
  1017 => x"2b527198",
  1018 => x"2ad40c71",
  1019 => x"902a7081",
  1020 => x"ff06d40c",
  1021 => x"5171882a",
  1022 => x"7081ff06",
  1023 => x"d40c5171",
  1024 => x"81ff06d4",
  1025 => x"0c72902a",
  1026 => x"7081ff06",
  1027 => x"d40c51d4",
  1028 => x"087081ff",
  1029 => x"06515182",
  1030 => x"b8bf5270",
  1031 => x"81ff2e09",
  1032 => x"81069438",
  1033 => x"81ff0bd4",
  1034 => x"0cd40870",
  1035 => x"81ff06ff",
  1036 => x"14545151",
  1037 => x"71e53870",
  1038 => x"bcd80c02",
  1039 => x"8c050d04",
  1040 => x"02fc050d",
  1041 => x"81c75181",
  1042 => x"ff0bd40c",
  1043 => x"ff115170",
  1044 => x"8025f438",
  1045 => x"0284050d",
  1046 => x"0402f005",
  1047 => x"0da0c02d",
  1048 => x"8fcf5380",
  1049 => x"5287fc80",
  1050 => x"f7519fce",
  1051 => x"2dbcd808",
  1052 => x"54bcd808",
  1053 => x"812e0981",
  1054 => x"06a33881",
  1055 => x"ff0bd40c",
  1056 => x"820a5284",
  1057 => x"9c80e951",
  1058 => x"9fce2dbc",
  1059 => x"d8088b38",
  1060 => x"81ff0bd4",
  1061 => x"0c7353a1",
  1062 => x"a304a0c0",
  1063 => x"2dff1353",
  1064 => x"72c13872",
  1065 => x"bcd80c02",
  1066 => x"90050d04",
  1067 => x"02f4050d",
  1068 => x"81ff0bd4",
  1069 => x"0c935380",
  1070 => x"5287fc80",
  1071 => x"c1519fce",
  1072 => x"2dbcd808",
  1073 => x"8b3881ff",
  1074 => x"0bd40c81",
  1075 => x"53a1d904",
  1076 => x"a0c02dff",
  1077 => x"135372df",
  1078 => x"3872bcd8",
  1079 => x"0c028c05",
  1080 => x"0d0402f0",
  1081 => x"050da0c0",
  1082 => x"2d83aa52",
  1083 => x"849c80c8",
  1084 => x"519fce2d",
  1085 => x"bcd80881",
  1086 => x"2e098106",
  1087 => x"92389f80",
  1088 => x"2dbcd808",
  1089 => x"83ffff06",
  1090 => x"537283aa",
  1091 => x"2e9738a1",
  1092 => x"ac2da2a0",
  1093 => x"048154a3",
  1094 => x"8504b98c",
  1095 => x"5185f22d",
  1096 => x"8054a385",
  1097 => x"0481ff0b",
  1098 => x"d40cb153",
  1099 => x"a0d92dbc",
  1100 => x"d808802e",
  1101 => x"80c03880",
  1102 => x"5287fc80",
  1103 => x"fa519fce",
  1104 => x"2dbcd808",
  1105 => x"b13881ff",
  1106 => x"0bd40cd4",
  1107 => x"085381ff",
  1108 => x"0bd40c81",
  1109 => x"ff0bd40c",
  1110 => x"81ff0bd4",
  1111 => x"0c81ff0b",
  1112 => x"d40c7286",
  1113 => x"2a708106",
  1114 => x"bcd80856",
  1115 => x"51537280",
  1116 => x"2e9338a2",
  1117 => x"95047282",
  1118 => x"2eff9f38",
  1119 => x"ff135372",
  1120 => x"ffaa3872",
  1121 => x"5473bcd8",
  1122 => x"0c029005",
  1123 => x"0d0402f0",
  1124 => x"050d810b",
  1125 => x"80c6cc0c",
  1126 => x"8454d008",
  1127 => x"708f2a70",
  1128 => x"81065151",
  1129 => x"5372f338",
  1130 => x"72d00ca0",
  1131 => x"c02db99c",
  1132 => x"5185f22d",
  1133 => x"d008708f",
  1134 => x"2a708106",
  1135 => x"51515372",
  1136 => x"f338810b",
  1137 => x"d00cb153",
  1138 => x"805284d4",
  1139 => x"80c0519f",
  1140 => x"ce2dbcd8",
  1141 => x"08812ea1",
  1142 => x"3872822e",
  1143 => x"0981068c",
  1144 => x"38b9a851",
  1145 => x"85f22d80",
  1146 => x"53a4af04",
  1147 => x"ff135372",
  1148 => x"d738ff14",
  1149 => x"5473ffa2",
  1150 => x"38a1e22d",
  1151 => x"bcd80880",
  1152 => x"c6cc0cbc",
  1153 => x"d8088b38",
  1154 => x"815287fc",
  1155 => x"80d0519f",
  1156 => x"ce2d81ff",
  1157 => x"0bd40cd0",
  1158 => x"08708f2a",
  1159 => x"70810651",
  1160 => x"515372f3",
  1161 => x"3872d00c",
  1162 => x"81ff0bd4",
  1163 => x"0c815372",
  1164 => x"bcd80c02",
  1165 => x"90050d04",
  1166 => x"02e8050d",
  1167 => x"785681ff",
  1168 => x"0bd40cd0",
  1169 => x"08708f2a",
  1170 => x"70810651",
  1171 => x"515372f3",
  1172 => x"3882810b",
  1173 => x"d00c81ff",
  1174 => x"0bd40c77",
  1175 => x"5287fc80",
  1176 => x"d8519fce",
  1177 => x"2dbcd808",
  1178 => x"802e8c38",
  1179 => x"b9c05185",
  1180 => x"f22d8153",
  1181 => x"a5ef0481",
  1182 => x"ff0bd40c",
  1183 => x"81fe0bd4",
  1184 => x"0c80ff55",
  1185 => x"75708405",
  1186 => x"57087098",
  1187 => x"2ad40c70",
  1188 => x"902c7081",
  1189 => x"ff06d40c",
  1190 => x"5470882c",
  1191 => x"7081ff06",
  1192 => x"d40c5470",
  1193 => x"81ff06d4",
  1194 => x"0c54ff15",
  1195 => x"55748025",
  1196 => x"d33881ff",
  1197 => x"0bd40c81",
  1198 => x"ff0bd40c",
  1199 => x"81ff0bd4",
  1200 => x"0c868da0",
  1201 => x"5481ff0b",
  1202 => x"d40cd408",
  1203 => x"81ff0655",
  1204 => x"748738ff",
  1205 => x"145473ed",
  1206 => x"3881ff0b",
  1207 => x"d40cd008",
  1208 => x"708f2a70",
  1209 => x"81065151",
  1210 => x"5372f338",
  1211 => x"72d00c72",
  1212 => x"bcd80c02",
  1213 => x"98050d04",
  1214 => x"02e8050d",
  1215 => x"78558056",
  1216 => x"81ff0bd4",
  1217 => x"0cd00870",
  1218 => x"8f2a7081",
  1219 => x"06515153",
  1220 => x"72f33882",
  1221 => x"810bd00c",
  1222 => x"81ff0bd4",
  1223 => x"0c775287",
  1224 => x"fc80d151",
  1225 => x"9fce2d80",
  1226 => x"dbc6df54",
  1227 => x"bcd80880",
  1228 => x"2e8a38b9",
  1229 => x"d05185f2",
  1230 => x"2da78f04",
  1231 => x"81ff0bd4",
  1232 => x"0cd40870",
  1233 => x"81ff0651",
  1234 => x"537281fe",
  1235 => x"2e098106",
  1236 => x"9d3880ff",
  1237 => x"539f802d",
  1238 => x"bcd80875",
  1239 => x"70840557",
  1240 => x"0cff1353",
  1241 => x"728025ed",
  1242 => x"388156a6",
  1243 => x"f404ff14",
  1244 => x"5473c938",
  1245 => x"81ff0bd4",
  1246 => x"0c81ff0b",
  1247 => x"d40cd008",
  1248 => x"708f2a70",
  1249 => x"81065151",
  1250 => x"5372f338",
  1251 => x"72d00c75",
  1252 => x"bcd80c02",
  1253 => x"98050d04",
  1254 => x"02f4050d",
  1255 => x"7470882a",
  1256 => x"83fe8006",
  1257 => x"7072982a",
  1258 => x"0772882b",
  1259 => x"87fc8080",
  1260 => x"0673982b",
  1261 => x"81f00a06",
  1262 => x"71730707",
  1263 => x"bcd80c56",
  1264 => x"51535102",
  1265 => x"8c050d04",
  1266 => x"02f8050d",
  1267 => x"028e0580",
  1268 => x"f52d7488",
  1269 => x"2b077083",
  1270 => x"ffff06bc",
  1271 => x"d80c5102",
  1272 => x"88050d04",
  1273 => x"02fc050d",
  1274 => x"72518071",
  1275 => x"0c800b84",
  1276 => x"120c0284",
  1277 => x"050d0402",
  1278 => x"f0050d75",
  1279 => x"70088412",
  1280 => x"08535353",
  1281 => x"ff547171",
  1282 => x"2ea838ab",
  1283 => x"bb2d8413",
  1284 => x"08708429",
  1285 => x"14881170",
  1286 => x"087081ff",
  1287 => x"06841808",
  1288 => x"81118706",
  1289 => x"841a0c53",
  1290 => x"51555151",
  1291 => x"51abb52d",
  1292 => x"715473bc",
  1293 => x"d80c0290",
  1294 => x"050d0402",
  1295 => x"f8050dab",
  1296 => x"bb2de008",
  1297 => x"708b2a70",
  1298 => x"81065152",
  1299 => x"5270802e",
  1300 => x"a13880c6",
  1301 => x"d0087084",
  1302 => x"2980c6d8",
  1303 => x"057381ff",
  1304 => x"06710c51",
  1305 => x"5180c6d0",
  1306 => x"08811187",
  1307 => x"0680c6d0",
  1308 => x"0c51800b",
  1309 => x"80c6f80c",
  1310 => x"abae2dab",
  1311 => x"b52d0288",
  1312 => x"050d0402",
  1313 => x"fc050dab",
  1314 => x"bb2d810b",
  1315 => x"80c6f80c",
  1316 => x"abb52d80",
  1317 => x"c6f80851",
  1318 => x"70f93802",
  1319 => x"84050d04",
  1320 => x"02fc050d",
  1321 => x"80c6d051",
  1322 => x"a7e42da8",
  1323 => x"bb51abaa",
  1324 => x"2daad42d",
  1325 => x"0284050d",
  1326 => x"0402f405",
  1327 => x"0daabb04",
  1328 => x"bcd80881",
  1329 => x"f02e0981",
  1330 => x"06893881",
  1331 => x"0bbccc0c",
  1332 => x"aabb04bc",
  1333 => x"d80881e0",
  1334 => x"2e098106",
  1335 => x"8938810b",
  1336 => x"bcd00caa",
  1337 => x"bb04bcd8",
  1338 => x"0852bcd0",
  1339 => x"08802e88",
  1340 => x"38bcd808",
  1341 => x"81800552",
  1342 => x"71842c72",
  1343 => x"8f065353",
  1344 => x"bccc0880",
  1345 => x"2e993872",
  1346 => x"8429bc8c",
  1347 => x"05721381",
  1348 => x"712b7009",
  1349 => x"73080673",
  1350 => x"0c515353",
  1351 => x"aab10472",
  1352 => x"8429bc8c",
  1353 => x"05721383",
  1354 => x"712b7208",
  1355 => x"07720c53",
  1356 => x"53800bbc",
  1357 => x"d00c800b",
  1358 => x"bccc0c80",
  1359 => x"c6d051a7",
  1360 => x"f72dbcd8",
  1361 => x"08ff24fe",
  1362 => x"f738800b",
  1363 => x"bcd80c02",
  1364 => x"8c050d04",
  1365 => x"02f8050d",
  1366 => x"bc8c528f",
  1367 => x"51807270",
  1368 => x"8405540c",
  1369 => x"ff115170",
  1370 => x"8025f238",
  1371 => x"0288050d",
  1372 => x"0402f005",
  1373 => x"0d7551ab",
  1374 => x"bb2d7082",
  1375 => x"2cfc06bc",
  1376 => x"8c117210",
  1377 => x"9e067108",
  1378 => x"70722a70",
  1379 => x"83068274",
  1380 => x"2b700974",
  1381 => x"06760c54",
  1382 => x"51565753",
  1383 => x"5153abb5",
  1384 => x"2d71bcd8",
  1385 => x"0c029005",
  1386 => x"0d047198",
  1387 => x"0c04ffb0",
  1388 => x"08bcd80c",
  1389 => x"04810bff",
  1390 => x"b00c0480",
  1391 => x"0bffb00c",
  1392 => x"0402fc05",
  1393 => x"0d810bbc",
  1394 => x"d40c8151",
  1395 => x"84e62d02",
  1396 => x"84050d04",
  1397 => x"02fc050d",
  1398 => x"800bbcd4",
  1399 => x"0c805184",
  1400 => x"e62d0284",
  1401 => x"050d0402",
  1402 => x"ec050d76",
  1403 => x"54805287",
  1404 => x"0b881580",
  1405 => x"f52d5653",
  1406 => x"74722483",
  1407 => x"38a05372",
  1408 => x"5182ef2d",
  1409 => x"81128b15",
  1410 => x"80f52d54",
  1411 => x"52727225",
  1412 => x"de380294",
  1413 => x"050d0402",
  1414 => x"f0050d80",
  1415 => x"c7880854",
  1416 => x"81f82d80",
  1417 => x"0b80c78c",
  1418 => x"0c730880",
  1419 => x"2e818438",
  1420 => x"820bbcec",
  1421 => x"0c80c78c",
  1422 => x"088f06bc",
  1423 => x"e80c7308",
  1424 => x"5271832e",
  1425 => x"96387183",
  1426 => x"26893871",
  1427 => x"812eaf38",
  1428 => x"ad9c0471",
  1429 => x"852e9f38",
  1430 => x"ad9c0488",
  1431 => x"1480f52d",
  1432 => x"841508b9",
  1433 => x"e0535452",
  1434 => x"85f22d71",
  1435 => x"84291370",
  1436 => x"085252ad",
  1437 => x"a0047351",
  1438 => x"abe72dad",
  1439 => x"9c0480c6",
  1440 => x"fc088815",
  1441 => x"082c7081",
  1442 => x"06515271",
  1443 => x"802e8738",
  1444 => x"b9e451ad",
  1445 => x"9904b9e8",
  1446 => x"5185f22d",
  1447 => x"84140851",
  1448 => x"85f22d80",
  1449 => x"c78c0881",
  1450 => x"0580c78c",
  1451 => x"0c8c1454",
  1452 => x"aca90402",
  1453 => x"90050d04",
  1454 => x"7180c788",
  1455 => x"0cac972d",
  1456 => x"80c78c08",
  1457 => x"ff0580c7",
  1458 => x"900c0402",
  1459 => x"e8050d80",
  1460 => x"c7880880",
  1461 => x"c7940857",
  1462 => x"5580f851",
  1463 => x"aaf12dbc",
  1464 => x"d808812a",
  1465 => x"70810651",
  1466 => x"52719b38",
  1467 => x"8751aaf1",
  1468 => x"2dbcd808",
  1469 => x"812a7081",
  1470 => x"06515271",
  1471 => x"802eb138",
  1472 => x"ae8604a9",
  1473 => x"b92d8751",
  1474 => x"aaf12dbc",
  1475 => x"d808f438",
  1476 => x"ae9604a9",
  1477 => x"b92d80f8",
  1478 => x"51aaf12d",
  1479 => x"bcd808f3",
  1480 => x"38bcd408",
  1481 => x"813270bc",
  1482 => x"d40c7052",
  1483 => x"5284e62d",
  1484 => x"800b80c7",
  1485 => x"800c800b",
  1486 => x"80c7840c",
  1487 => x"bcd40882",
  1488 => x"fd3880da",
  1489 => x"51aaf12d",
  1490 => x"bcd80880",
  1491 => x"2e8c3880",
  1492 => x"c7800881",
  1493 => x"800780c7",
  1494 => x"800c80d9",
  1495 => x"51aaf12d",
  1496 => x"bcd80880",
  1497 => x"2e8c3880",
  1498 => x"c7800880",
  1499 => x"c00780c7",
  1500 => x"800c8194",
  1501 => x"51aaf12d",
  1502 => x"bcd80880",
  1503 => x"2e8b3880",
  1504 => x"c7800890",
  1505 => x"0780c780",
  1506 => x"0c819151",
  1507 => x"aaf12dbc",
  1508 => x"d808802e",
  1509 => x"8b3880c7",
  1510 => x"8008a007",
  1511 => x"80c7800c",
  1512 => x"81f551aa",
  1513 => x"f12dbcd8",
  1514 => x"08802e8b",
  1515 => x"3880c780",
  1516 => x"08810780",
  1517 => x"c7800c81",
  1518 => x"f251aaf1",
  1519 => x"2dbcd808",
  1520 => x"802e8b38",
  1521 => x"80c78008",
  1522 => x"820780c7",
  1523 => x"800c81eb",
  1524 => x"51aaf12d",
  1525 => x"bcd80880",
  1526 => x"2e8b3880",
  1527 => x"c7800884",
  1528 => x"0780c780",
  1529 => x"0c81f451",
  1530 => x"aaf12dbc",
  1531 => x"d808802e",
  1532 => x"8b3880c7",
  1533 => x"80088807",
  1534 => x"80c7800c",
  1535 => x"80d851aa",
  1536 => x"f12dbcd8",
  1537 => x"08802e8c",
  1538 => x"3880c784",
  1539 => x"08818007",
  1540 => x"80c7840c",
  1541 => x"9251aaf1",
  1542 => x"2dbcd808",
  1543 => x"802e8c38",
  1544 => x"80c78408",
  1545 => x"80c00780",
  1546 => x"c7840c94",
  1547 => x"51aaf12d",
  1548 => x"bcd80880",
  1549 => x"2e8b3880",
  1550 => x"c7840890",
  1551 => x"0780c784",
  1552 => x"0c9151aa",
  1553 => x"f12dbcd8",
  1554 => x"08802e8b",
  1555 => x"3880c784",
  1556 => x"08a00780",
  1557 => x"c7840c9d",
  1558 => x"51aaf12d",
  1559 => x"bcd80880",
  1560 => x"2e8b3880",
  1561 => x"c7840881",
  1562 => x"0780c784",
  1563 => x"0c9b51aa",
  1564 => x"f12dbcd8",
  1565 => x"08802e8b",
  1566 => x"3880c784",
  1567 => x"08820780",
  1568 => x"c7840c9c",
  1569 => x"51aaf12d",
  1570 => x"bcd80880",
  1571 => x"2e8b3880",
  1572 => x"c7840884",
  1573 => x"0780c784",
  1574 => x"0ca351aa",
  1575 => x"f12dbcd8",
  1576 => x"08802e8b",
  1577 => x"3880c784",
  1578 => x"08880780",
  1579 => x"c7840c81",
  1580 => x"fd51aaf1",
  1581 => x"2d81fa51",
  1582 => x"aaf12db7",
  1583 => x"860481f5",
  1584 => x"51aaf12d",
  1585 => x"bcd80881",
  1586 => x"2a708106",
  1587 => x"51527180",
  1588 => x"2eb33880",
  1589 => x"c7900852",
  1590 => x"71802e8a",
  1591 => x"38ff1280",
  1592 => x"c7900cb2",
  1593 => x"850480c7",
  1594 => x"8c081080",
  1595 => x"c78c0805",
  1596 => x"70842916",
  1597 => x"51528812",
  1598 => x"08802e89",
  1599 => x"38ff5188",
  1600 => x"12085271",
  1601 => x"2d81f251",
  1602 => x"aaf12dbc",
  1603 => x"d808812a",
  1604 => x"70810651",
  1605 => x"5271802e",
  1606 => x"b43880c7",
  1607 => x"8c08ff11",
  1608 => x"80c79008",
  1609 => x"56535373",
  1610 => x"72258a38",
  1611 => x"811480c7",
  1612 => x"900cb2cd",
  1613 => x"04721013",
  1614 => x"70842916",
  1615 => x"51528812",
  1616 => x"08802e89",
  1617 => x"38fe5188",
  1618 => x"12085271",
  1619 => x"2d81fd51",
  1620 => x"aaf12dbc",
  1621 => x"d808812a",
  1622 => x"70810651",
  1623 => x"5271802e",
  1624 => x"b13880c7",
  1625 => x"9008802e",
  1626 => x"8a38800b",
  1627 => x"80c7900c",
  1628 => x"b3920480",
  1629 => x"c78c0810",
  1630 => x"80c78c08",
  1631 => x"05708429",
  1632 => x"16515288",
  1633 => x"1208802e",
  1634 => x"8938fd51",
  1635 => x"88120852",
  1636 => x"712d81fa",
  1637 => x"51aaf12d",
  1638 => x"bcd80881",
  1639 => x"2a708106",
  1640 => x"51527180",
  1641 => x"2eb13880",
  1642 => x"c78c08ff",
  1643 => x"11545280",
  1644 => x"c7900873",
  1645 => x"25893872",
  1646 => x"80c7900c",
  1647 => x"b3d70471",
  1648 => x"10127084",
  1649 => x"29165152",
  1650 => x"88120880",
  1651 => x"2e8938fc",
  1652 => x"51881208",
  1653 => x"52712d80",
  1654 => x"c7900870",
  1655 => x"53547380",
  1656 => x"2e8a388c",
  1657 => x"15ff1555",
  1658 => x"55b3de04",
  1659 => x"820bbcec",
  1660 => x"0c718f06",
  1661 => x"bce80c81",
  1662 => x"eb51aaf1",
  1663 => x"2dbcd808",
  1664 => x"812a7081",
  1665 => x"06515271",
  1666 => x"802ead38",
  1667 => x"7408852e",
  1668 => x"098106a4",
  1669 => x"38881580",
  1670 => x"f52dff05",
  1671 => x"52718816",
  1672 => x"81b72d71",
  1673 => x"982b5271",
  1674 => x"80258838",
  1675 => x"800b8816",
  1676 => x"81b72d74",
  1677 => x"51abe72d",
  1678 => x"81f451aa",
  1679 => x"f12dbcd8",
  1680 => x"08812a70",
  1681 => x"81065152",
  1682 => x"71802eb3",
  1683 => x"38740885",
  1684 => x"2e098106",
  1685 => x"aa388815",
  1686 => x"80f52d81",
  1687 => x"05527188",
  1688 => x"1681b72d",
  1689 => x"7181ff06",
  1690 => x"8b1680f5",
  1691 => x"2d545272",
  1692 => x"72278738",
  1693 => x"72881681",
  1694 => x"b72d7451",
  1695 => x"abe72d80",
  1696 => x"da51aaf1",
  1697 => x"2dbcd808",
  1698 => x"812a7081",
  1699 => x"06515271",
  1700 => x"802e81ac",
  1701 => x"3880c788",
  1702 => x"0880c790",
  1703 => x"08555373",
  1704 => x"802e8a38",
  1705 => x"8c13ff15",
  1706 => x"5553b59f",
  1707 => x"04720852",
  1708 => x"71822ea6",
  1709 => x"38718226",
  1710 => x"89387181",
  1711 => x"2eaa38b6",
  1712 => x"c0047183",
  1713 => x"2eb43871",
  1714 => x"842e0981",
  1715 => x"0680f138",
  1716 => x"88130851",
  1717 => x"adb82db6",
  1718 => x"c00480c7",
  1719 => x"90085188",
  1720 => x"13085271",
  1721 => x"2db6c004",
  1722 => x"810b8814",
  1723 => x"082b80c6",
  1724 => x"fc083280",
  1725 => x"c6fc0cb6",
  1726 => x"95048813",
  1727 => x"80f52d81",
  1728 => x"058b1480",
  1729 => x"f52d5354",
  1730 => x"71742483",
  1731 => x"38805473",
  1732 => x"881481b7",
  1733 => x"2dac972d",
  1734 => x"b6c00475",
  1735 => x"08802ea3",
  1736 => x"38750851",
  1737 => x"aaf12dbc",
  1738 => x"d8088106",
  1739 => x"5271802e",
  1740 => x"8c3880c7",
  1741 => x"90085184",
  1742 => x"16085271",
  1743 => x"2d881656",
  1744 => x"75d93880",
  1745 => x"54800bbc",
  1746 => x"ec0c738f",
  1747 => x"06bce80c",
  1748 => x"a0527380",
  1749 => x"c790082e",
  1750 => x"09810699",
  1751 => x"3880c78c",
  1752 => x"08ff0574",
  1753 => x"32700981",
  1754 => x"05707207",
  1755 => x"9f2a9171",
  1756 => x"31515153",
  1757 => x"53715182",
  1758 => x"ef2d8114",
  1759 => x"548e7425",
  1760 => x"c438bcd4",
  1761 => x"085271bc",
  1762 => x"d80c0298",
  1763 => x"050d0400",
  1764 => x"00ffffff",
  1765 => x"ff00ffff",
  1766 => x"ffff00ff",
  1767 => x"ffffff00",
  1768 => x"52657365",
  1769 => x"74000000",
  1770 => x"53617665",
  1771 => x"20736574",
  1772 => x"74696e67",
  1773 => x"73000000",
  1774 => x"5363616e",
  1775 => x"6c696e65",
  1776 => x"73000000",
  1777 => x"4c6f6164",
  1778 => x"20524f4d",
  1779 => x"20100000",
  1780 => x"45786974",
  1781 => x"00000000",
  1782 => x"56474120",
  1783 => x"2d203331",
  1784 => x"4b487a2c",
  1785 => x"20363048",
  1786 => x"7a000000",
  1787 => x"5456202d",
  1788 => x"20343830",
  1789 => x"692c2036",
  1790 => x"30487a00",
  1791 => x"4261636b",
  1792 => x"00000000",
  1793 => x"46504741",
  1794 => x"47454e20",
  1795 => x"43464700",
  1796 => x"496e6974",
  1797 => x"69616c69",
  1798 => x"7a696e67",
  1799 => x"20534420",
  1800 => x"63617264",
  1801 => x"0a000000",
  1802 => x"424f4f54",
  1803 => x"20202020",
  1804 => x"47454e00",
  1805 => x"43617264",
  1806 => x"20696e69",
  1807 => x"74206661",
  1808 => x"696c6564",
  1809 => x"0a000000",
  1810 => x"4d425220",
  1811 => x"6661696c",
  1812 => x"0a000000",
  1813 => x"46415431",
  1814 => x"36202020",
  1815 => x"00000000",
  1816 => x"46415433",
  1817 => x"32202020",
  1818 => x"00000000",
  1819 => x"4e6f2070",
  1820 => x"61727469",
  1821 => x"74696f6e",
  1822 => x"20736967",
  1823 => x"0a000000",
  1824 => x"42616420",
  1825 => x"70617274",
  1826 => x"0a000000",
  1827 => x"53444843",
  1828 => x"20657272",
  1829 => x"6f72210a",
  1830 => x"00000000",
  1831 => x"53442069",
  1832 => x"6e69742e",
  1833 => x"2e2e0a00",
  1834 => x"53442063",
  1835 => x"61726420",
  1836 => x"72657365",
  1837 => x"74206661",
  1838 => x"696c6564",
  1839 => x"210a0000",
  1840 => x"57726974",
  1841 => x"65206661",
  1842 => x"696c6564",
  1843 => x"0a000000",
  1844 => x"52656164",
  1845 => x"20666169",
  1846 => x"6c65640a",
  1847 => x"00000000",
  1848 => x"16200000",
  1849 => x"14200000",
  1850 => x"15200000",
  1851 => x"00000002",
  1852 => x"00000000",
  1853 => x"00000002",
  1854 => x"00001ba0",
  1855 => x"0000049a",
  1856 => x"00000002",
  1857 => x"00001ba8",
  1858 => x"0000036d",
  1859 => x"00000003",
  1860 => x"00001d48",
  1861 => x"00000002",
  1862 => x"00000001",
  1863 => x"00001bb8",
  1864 => x"00000001",
  1865 => x"00000002",
  1866 => x"00001bc4",
  1867 => x"00000734",
  1868 => x"00000002",
  1869 => x"00001bd0",
  1870 => x"000015d4",
  1871 => x"00000000",
  1872 => x"00000000",
  1873 => x"00000000",
  1874 => x"00001bd8",
  1875 => x"00001bec",
  1876 => x"00000002",
  1877 => x"00001e88",
  1878 => x"00000528",
  1879 => x"00000002",
  1880 => x"00001ea6",
  1881 => x"00000528",
  1882 => x"00000002",
  1883 => x"00001ec4",
  1884 => x"00000528",
  1885 => x"00000002",
  1886 => x"00001ee2",
  1887 => x"00000528",
  1888 => x"00000002",
  1889 => x"00001f00",
  1890 => x"00000528",
  1891 => x"00000002",
  1892 => x"00001f1e",
  1893 => x"00000528",
  1894 => x"00000002",
  1895 => x"00001f3c",
  1896 => x"00000528",
  1897 => x"00000002",
  1898 => x"00001f5a",
  1899 => x"00000528",
  1900 => x"00000002",
  1901 => x"00001f78",
  1902 => x"00000528",
  1903 => x"00000002",
  1904 => x"00001f96",
  1905 => x"00000528",
  1906 => x"00000002",
  1907 => x"00001fb4",
  1908 => x"00000528",
  1909 => x"00000002",
  1910 => x"00001fd2",
  1911 => x"00000528",
  1912 => x"00000002",
  1913 => x"00001ff0",
  1914 => x"00000528",
  1915 => x"00000004",
  1916 => x"00001bfc",
  1917 => x"00001cf4",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"000006c8",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"00000000",
  1932 => x"00000000",
  1933 => x"00000000",
  1934 => x"00000000",
  1935 => x"00000000",
  1936 => x"00000000",
  1937 => x"00000000",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

