-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbc",
     9 => x"8c080b0b",
    10 => x"0bbc9008",
    11 => x"0b0b0bbc",
    12 => x"94080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bc940c0b",
    16 => x"0b0bbc90",
    17 => x"0c0b0b0b",
    18 => x"bc8c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb6c8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bc8c7080",
    57 => x"c6cc278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518edf04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbc9c0c",
    65 => x"9f0bbca0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bca008ff",
    69 => x"05bca00c",
    70 => x"bca00880",
    71 => x"25eb38bc",
    72 => x"9c08ff05",
    73 => x"bc9c0cbc",
    74 => x"9c088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbc",
    94 => x"9c08258f",
    95 => x"3882b32d",
    96 => x"bc9c08ff",
    97 => x"05bc9c0c",
    98 => x"82f504bc",
    99 => x"9c08bca0",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038bc9c",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"bca00881",
   109 => x"05bca00c",
   110 => x"bca00851",
   111 => x"9f7125e2",
   112 => x"38800bbc",
   113 => x"a00cbc9c",
   114 => x"088105bc",
   115 => x"9c0c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34bca008",
   120 => x"8105bca0",
   121 => x"0cbca008",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbca00c",
   125 => x"bc9c0881",
   126 => x"05bc9c0c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"bca40cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbc",
   162 => x"a40c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72bca408",
   167 => x"8407bca4",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"b9a40c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"bca40852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"fc050d72",
   198 => x"70820680",
   199 => x"c6b00c70",
   200 => x"81065151",
   201 => x"70b9c80b",
   202 => x"81b72d70",
   203 => x"bc8c0c02",
   204 => x"84050d04",
   205 => x"02f8050d",
   206 => x"b7bc52bc",
   207 => x"a8519ba6",
   208 => x"2dbc8c08",
   209 => x"802e9d38",
   210 => x"bfc452bc",
   211 => x"a8519de5",
   212 => x"2dbfc408",
   213 => x"bcb40cbf",
   214 => x"c408fec0",
   215 => x"0cbfc408",
   216 => x"5186932d",
   217 => x"0288050d",
   218 => x"0402f005",
   219 => x"0d805191",
   220 => x"912db7bc",
   221 => x"52bca851",
   222 => x"9ba62dbc",
   223 => x"8c08802e",
   224 => x"a538bcb4",
   225 => x"08bfc40c",
   226 => x"bfc85480",
   227 => x"fd538074",
   228 => x"70840556",
   229 => x"0cff1353",
   230 => x"728025f2",
   231 => x"38bfc452",
   232 => x"bca8519e",
   233 => x"8e2d0290",
   234 => x"050d0402",
   235 => x"d8050dbc",
   236 => x"b408fec0",
   237 => x"0c810bfe",
   238 => x"c40c840b",
   239 => x"fec40c7b",
   240 => x"52bca851",
   241 => x"9ba62dbc",
   242 => x"8c0853bc",
   243 => x"8c08802e",
   244 => x"81a438bc",
   245 => x"ac085580",
   246 => x"0bff1657",
   247 => x"5975792e",
   248 => x"8b388119",
   249 => x"76812a57",
   250 => x"5975f738",
   251 => x"f7195974",
   252 => x"b080802e",
   253 => x"09810689",
   254 => x"38820bfe",
   255 => x"dc0c8898",
   256 => x"04749880",
   257 => x"802e0981",
   258 => x"06893881",
   259 => x"0bfedc0c",
   260 => x"88980480",
   261 => x"0bfedc0c",
   262 => x"815a8075",
   263 => x"2580d538",
   264 => x"78527551",
   265 => x"84812dbf",
   266 => x"c452bca8",
   267 => x"519de52d",
   268 => x"bc8c0880",
   269 => x"2ea738bf",
   270 => x"c45883fc",
   271 => x"57777084",
   272 => x"05590870",
   273 => x"83ffff06",
   274 => x"71902afe",
   275 => x"c80cfec8",
   276 => x"0cfc1858",
   277 => x"53768025",
   278 => x"e43888e4",
   279 => x"04bc8c08",
   280 => x"5a848055",
   281 => x"bca8519d",
   282 => x"b72dfc80",
   283 => x"15811757",
   284 => x"55889a04",
   285 => x"795372bc",
   286 => x"8c0c02a8",
   287 => x"050d0402",
   288 => x"fc050dab",
   289 => x"8b2dfec4",
   290 => x"5181710c",
   291 => x"82710c02",
   292 => x"84050d04",
   293 => x"02f4050d",
   294 => x"74767853",
   295 => x"54528071",
   296 => x"25973872",
   297 => x"70810554",
   298 => x"80f52d72",
   299 => x"70810554",
   300 => x"81b72dff",
   301 => x"115170eb",
   302 => x"38807281",
   303 => x"b72d028c",
   304 => x"050d0402",
   305 => x"e8050d77",
   306 => x"56807056",
   307 => x"54737624",
   308 => x"b33880c5",
   309 => x"d408742e",
   310 => x"ab387351",
   311 => x"98f12dbc",
   312 => x"8c08bc8c",
   313 => x"08098105",
   314 => x"70bc8c08",
   315 => x"079f2a77",
   316 => x"05811757",
   317 => x"57535374",
   318 => x"76248938",
   319 => x"80c5d408",
   320 => x"7426d738",
   321 => x"72bc8c0c",
   322 => x"0298050d",
   323 => x"0402f405",
   324 => x"0dbbb808",
   325 => x"155189c3",
   326 => x"2dbc8c08",
   327 => x"802e9538",
   328 => x"8b53bc8c",
   329 => x"085280c3",
   330 => x"c4518994",
   331 => x"2d80c3c4",
   332 => x"5187ab2d",
   333 => x"b9a851ac",
   334 => x"ef2dab8b",
   335 => x"2d805184",
   336 => x"e62d028c",
   337 => x"050d0402",
   338 => x"dc050d80",
   339 => x"705a5574",
   340 => x"bbb80825",
   341 => x"b13880c5",
   342 => x"d408752e",
   343 => x"a9387851",
   344 => x"98f12dbc",
   345 => x"8c080981",
   346 => x"0570bc8c",
   347 => x"08079f2a",
   348 => x"7605811b",
   349 => x"5b565474",
   350 => x"bbb80825",
   351 => x"893880c5",
   352 => x"d4087926",
   353 => x"d9388055",
   354 => x"7880c5d4",
   355 => x"082781d0",
   356 => x"38785198",
   357 => x"f12dbc8c",
   358 => x"08802e81",
   359 => x"a538bc8c",
   360 => x"088b0580",
   361 => x"f52d7084",
   362 => x"2a708106",
   363 => x"77107884",
   364 => x"2b80c3c4",
   365 => x"0b80f52d",
   366 => x"5c5c5351",
   367 => x"55567380",
   368 => x"2e80c738",
   369 => x"7416822b",
   370 => x"8d830bba",
   371 => x"8c120c54",
   372 => x"77753110",
   373 => x"bcbc1155",
   374 => x"56907470",
   375 => x"81055681",
   376 => x"b72da074",
   377 => x"81b72d76",
   378 => x"81ff0681",
   379 => x"16585473",
   380 => x"802e8a38",
   381 => x"9c5380c3",
   382 => x"c4528c83",
   383 => x"048b53bc",
   384 => x"8c0852bc",
   385 => x"be16518c",
   386 => x"ba047416",
   387 => x"822b8a8d",
   388 => x"0bba8c12",
   389 => x"0c547681",
   390 => x"ff068116",
   391 => x"58547380",
   392 => x"2e8a389c",
   393 => x"5380c3c4",
   394 => x"528cb204",
   395 => x"8b53bc8c",
   396 => x"08527775",
   397 => x"3110bcbc",
   398 => x"05517655",
   399 => x"89942d8c",
   400 => x"d5047490",
   401 => x"29753170",
   402 => x"10bcbc05",
   403 => x"5154bc8c",
   404 => x"087481b7",
   405 => x"2d811959",
   406 => x"748b24a2",
   407 => x"388b8804",
   408 => x"74902975",
   409 => x"317010bc",
   410 => x"bc058c77",
   411 => x"31575154",
   412 => x"807481b7",
   413 => x"2d9e14ff",
   414 => x"16565474",
   415 => x"f33802a4",
   416 => x"050d0402",
   417 => x"fc050dbb",
   418 => x"b8081351",
   419 => x"89c32dbc",
   420 => x"8c08802e",
   421 => x"8838bc8c",
   422 => x"08519191",
   423 => x"2d800bbb",
   424 => x"b80c8ac7",
   425 => x"2dabce2d",
   426 => x"0284050d",
   427 => x"0402fc05",
   428 => x"0d725170",
   429 => x"fd2ead38",
   430 => x"70fd248a",
   431 => x"3870fc2e",
   432 => x"80c4388e",
   433 => x"8e0470fe",
   434 => x"2eb13870",
   435 => x"ff2e0981",
   436 => x"06bc38bb",
   437 => x"b8085170",
   438 => x"802eb338",
   439 => x"ff11bbb8",
   440 => x"0c8e8e04",
   441 => x"bbb808f0",
   442 => x"0570bbb8",
   443 => x"0c517080",
   444 => x"259c3880",
   445 => x"0bbbb80c",
   446 => x"8e8e04bb",
   447 => x"b8088105",
   448 => x"bbb80c8e",
   449 => x"8e04bbb8",
   450 => x"089005bb",
   451 => x"b80c8ac7",
   452 => x"2dabce2d",
   453 => x"0284050d",
   454 => x"0402fc05",
   455 => x"0d800bbb",
   456 => x"b80c8ac7",
   457 => x"2dba8451",
   458 => x"acef2d02",
   459 => x"84050d04",
   460 => x"02f8050d",
   461 => x"80c6b008",
   462 => x"8206b9c8",
   463 => x"0b80f52d",
   464 => x"52527080",
   465 => x"2e853871",
   466 => x"810752bc",
   467 => x"b808802e",
   468 => x"85387190",
   469 => x"075271bc",
   470 => x"8c0c0288",
   471 => x"050d0402",
   472 => x"f4050d81",
   473 => x"0bbcb80c",
   474 => x"90518693",
   475 => x"2d810bfe",
   476 => x"c40c860b",
   477 => x"fec40ca8",
   478 => x"d72daaec",
   479 => x"2da8ba2d",
   480 => x"a8ba2d81",
   481 => x"f82d8151",
   482 => x"84e62da8",
   483 => x"ba2da8ba",
   484 => x"2d815184",
   485 => x"e62d830b",
   486 => x"fecc0cb7",
   487 => x"c85185f2",
   488 => x"2d8452a2",
   489 => x"c52d92b2",
   490 => x"2dbc8c08",
   491 => x"802e8638",
   492 => x"fe528fbd",
   493 => x"04ff1252",
   494 => x"718024e7",
   495 => x"3871802e",
   496 => x"81813886",
   497 => x"b42db7e0",
   498 => x"5187ab2d",
   499 => x"bc8c0880",
   500 => x"2e8f38b9",
   501 => x"a851acef",
   502 => x"2d805184",
   503 => x"e62d8feb",
   504 => x"04bc8c08",
   505 => x"518e992d",
   506 => x"aaf82d82",
   507 => x"0bfec40c",
   508 => x"a8f02dad",
   509 => x"822dbc8c",
   510 => x"0880c6b4",
   511 => x"08882b80",
   512 => x"c6b80807",
   513 => x"fed80c53",
   514 => x"8eb02dbc",
   515 => x"8c08bcb4",
   516 => x"082ea238",
   517 => x"bc8c08bc",
   518 => x"b40cbc8c",
   519 => x"08fec00c",
   520 => x"84527251",
   521 => x"84e62da8",
   522 => x"ba2da8ba",
   523 => x"2dff1252",
   524 => x"718025ee",
   525 => x"3872802e",
   526 => x"ffb1388a",
   527 => x"0bfec40c",
   528 => x"8ff004b7",
   529 => x"ec5185f2",
   530 => x"2d800bbc",
   531 => x"8c0c028c",
   532 => x"050d0402",
   533 => x"e8050d77",
   534 => x"797b5855",
   535 => x"55805372",
   536 => x"7625a338",
   537 => x"74708105",
   538 => x"5680f52d",
   539 => x"74708105",
   540 => x"5680f52d",
   541 => x"52527171",
   542 => x"2e863881",
   543 => x"51918804",
   544 => x"81135390",
   545 => x"df048051",
   546 => x"70bc8c0c",
   547 => x"0298050d",
   548 => x"0402ec05",
   549 => x"0d765574",
   550 => x"802ebe38",
   551 => x"9a1580e0",
   552 => x"2d51a6ff",
   553 => x"2dbc8c08",
   554 => x"bc8c0880",
   555 => x"c5f40cbc",
   556 => x"8c085454",
   557 => x"80c5d008",
   558 => x"802e9938",
   559 => x"941580e0",
   560 => x"2d51a6ff",
   561 => x"2dbc8c08",
   562 => x"902b83ff",
   563 => x"f00a0670",
   564 => x"75075153",
   565 => x"7280c5f4",
   566 => x"0c80c5f4",
   567 => x"08537280",
   568 => x"2e9d3880",
   569 => x"c5c808fe",
   570 => x"14712980",
   571 => x"c5dc0805",
   572 => x"80c5f80c",
   573 => x"70842b80",
   574 => x"c5d40c54",
   575 => x"92ad0480",
   576 => x"c5e00880",
   577 => x"c5f40c80",
   578 => x"c5e40880",
   579 => x"c5f80c80",
   580 => x"c5d00880",
   581 => x"2e8b3880",
   582 => x"c5c80884",
   583 => x"2b5392a8",
   584 => x"0480c5e8",
   585 => x"08842b53",
   586 => x"7280c5d4",
   587 => x"0c029405",
   588 => x"0d0402d8",
   589 => x"050d800b",
   590 => x"80c5d00c",
   591 => x"bfc45280",
   592 => x"51a5af2d",
   593 => x"bc8c0854",
   594 => x"bc8c088c",
   595 => x"38b88051",
   596 => x"85f22d73",
   597 => x"5597f704",
   598 => x"8056810b",
   599 => x"80c5fc0c",
   600 => x"8853b88c",
   601 => x"52bffa51",
   602 => x"90d32dbc",
   603 => x"8c08762e",
   604 => x"09810688",
   605 => x"38bc8c08",
   606 => x"80c5fc0c",
   607 => x"8853b898",
   608 => x"5280c096",
   609 => x"5190d32d",
   610 => x"bc8c0888",
   611 => x"38bc8c08",
   612 => x"80c5fc0c",
   613 => x"80c5fc08",
   614 => x"802e80fc",
   615 => x"3880c38a",
   616 => x"0b80f52d",
   617 => x"80c38b0b",
   618 => x"80f52d71",
   619 => x"982b7190",
   620 => x"2b0780c3",
   621 => x"8c0b80f5",
   622 => x"2d70882b",
   623 => x"720780c3",
   624 => x"8d0b80f5",
   625 => x"2d710780",
   626 => x"c3c20b80",
   627 => x"f52d80c3",
   628 => x"c30b80f5",
   629 => x"2d71882b",
   630 => x"07535f54",
   631 => x"525a5657",
   632 => x"557381ab",
   633 => x"aa2e0981",
   634 => x"068d3875",
   635 => x"51a6cf2d",
   636 => x"bc8c0856",
   637 => x"94840473",
   638 => x"82d4d52e",
   639 => x"8738b8a4",
   640 => x"5194c704",
   641 => x"bfc45275",
   642 => x"51a5af2d",
   643 => x"bc8c0855",
   644 => x"bc8c0880",
   645 => x"2e83e038",
   646 => x"8853b898",
   647 => x"5280c096",
   648 => x"5190d32d",
   649 => x"bc8c088a",
   650 => x"38810b80",
   651 => x"c5d00c94",
   652 => x"cd048853",
   653 => x"b88c52bf",
   654 => x"fa5190d3",
   655 => x"2dbc8c08",
   656 => x"802e8a38",
   657 => x"b8b85185",
   658 => x"f22d95a9",
   659 => x"0480c3c2",
   660 => x"0b80f52d",
   661 => x"547380d5",
   662 => x"2e098106",
   663 => x"80cb3880",
   664 => x"c3c30b80",
   665 => x"f52d5473",
   666 => x"81aa2e09",
   667 => x"8106ba38",
   668 => x"800bbfc4",
   669 => x"0b80f52d",
   670 => x"56547481",
   671 => x"e92e8338",
   672 => x"81547481",
   673 => x"eb2e8c38",
   674 => x"80557375",
   675 => x"2e098106",
   676 => x"82e538bf",
   677 => x"cf0b80f5",
   678 => x"2d55748d",
   679 => x"38bfd00b",
   680 => x"80f52d54",
   681 => x"73822e86",
   682 => x"38805597",
   683 => x"f704bfd1",
   684 => x"0b80f52d",
   685 => x"7080c5c8",
   686 => x"0cff0580",
   687 => x"c5cc0cbf",
   688 => x"d20b80f5",
   689 => x"2dbfd30b",
   690 => x"80f52d58",
   691 => x"76057782",
   692 => x"80290570",
   693 => x"80c5d80c",
   694 => x"bfd40b80",
   695 => x"f52d7080",
   696 => x"c5ec0c80",
   697 => x"c5d00859",
   698 => x"57587680",
   699 => x"2e81ad38",
   700 => x"8853b898",
   701 => x"5280c096",
   702 => x"5190d32d",
   703 => x"bc8c0881",
   704 => x"f63880c5",
   705 => x"c8087084",
   706 => x"2b80c5d4",
   707 => x"0c7080c5",
   708 => x"e80cbfe9",
   709 => x"0b80f52d",
   710 => x"bfe80b80",
   711 => x"f52d7182",
   712 => x"802905bf",
   713 => x"ea0b80f5",
   714 => x"2d708480",
   715 => x"802912bf",
   716 => x"eb0b80f5",
   717 => x"2d708180",
   718 => x"0a291270",
   719 => x"80c5f00c",
   720 => x"80c5ec08",
   721 => x"712980c5",
   722 => x"d8080570",
   723 => x"80c5dc0c",
   724 => x"bff10b80",
   725 => x"f52dbff0",
   726 => x"0b80f52d",
   727 => x"71828029",
   728 => x"05bff20b",
   729 => x"80f52d70",
   730 => x"84808029",
   731 => x"12bff30b",
   732 => x"80f52d70",
   733 => x"982b81f0",
   734 => x"0a067205",
   735 => x"7080c5e0",
   736 => x"0cfe117e",
   737 => x"29770580",
   738 => x"c5e40c52",
   739 => x"59524354",
   740 => x"5e515259",
   741 => x"525d5759",
   742 => x"5797f004",
   743 => x"bfd60b80",
   744 => x"f52dbfd5",
   745 => x"0b80f52d",
   746 => x"71828029",
   747 => x"057080c5",
   748 => x"d40c70a0",
   749 => x"2983ff05",
   750 => x"70892a70",
   751 => x"80c5e80c",
   752 => x"bfdb0b80",
   753 => x"f52dbfda",
   754 => x"0b80f52d",
   755 => x"71828029",
   756 => x"057080c5",
   757 => x"f00c7b71",
   758 => x"291e7080",
   759 => x"c5e40c7d",
   760 => x"80c5e00c",
   761 => x"730580c5",
   762 => x"dc0c555e",
   763 => x"51515555",
   764 => x"80519191",
   765 => x"2d815574",
   766 => x"bc8c0c02",
   767 => x"a8050d04",
   768 => x"02ec050d",
   769 => x"7670872c",
   770 => x"7180ff06",
   771 => x"55565480",
   772 => x"c5d0088a",
   773 => x"3873882c",
   774 => x"7481ff06",
   775 => x"5455bfc4",
   776 => x"5280c5d8",
   777 => x"081551a5",
   778 => x"af2dbc8c",
   779 => x"0854bc8c",
   780 => x"08802eb4",
   781 => x"3880c5d0",
   782 => x"08802e98",
   783 => x"38728429",
   784 => x"bfc40570",
   785 => x"085253a6",
   786 => x"cf2dbc8c",
   787 => x"08f00a06",
   788 => x"5398e604",
   789 => x"7210bfc4",
   790 => x"057080e0",
   791 => x"2d5253a6",
   792 => x"ff2dbc8c",
   793 => x"08537254",
   794 => x"73bc8c0c",
   795 => x"0294050d",
   796 => x"0402e005",
   797 => x"0d797084",
   798 => x"2c80c5f8",
   799 => x"0805718f",
   800 => x"06525553",
   801 => x"728938bf",
   802 => x"c4527351",
   803 => x"a5af2d72",
   804 => x"a029bfc4",
   805 => x"05548074",
   806 => x"80f52d56",
   807 => x"5374732e",
   808 => x"83388153",
   809 => x"7481e52e",
   810 => x"81f13881",
   811 => x"70740654",
   812 => x"5872802e",
   813 => x"81e5388b",
   814 => x"1480f52d",
   815 => x"70832a79",
   816 => x"06585676",
   817 => x"9938bbbc",
   818 => x"08537289",
   819 => x"387280c3",
   820 => x"c40b81b7",
   821 => x"2d76bbbc",
   822 => x"0c73539b",
   823 => x"9d04758f",
   824 => x"2e098106",
   825 => x"81b53874",
   826 => x"9f068d29",
   827 => x"80c3b711",
   828 => x"51538114",
   829 => x"80f52d73",
   830 => x"70810555",
   831 => x"81b72d83",
   832 => x"1480f52d",
   833 => x"73708105",
   834 => x"5581b72d",
   835 => x"851480f5",
   836 => x"2d737081",
   837 => x"055581b7",
   838 => x"2d871480",
   839 => x"f52d7370",
   840 => x"81055581",
   841 => x"b72d8914",
   842 => x"80f52d73",
   843 => x"70810555",
   844 => x"81b72d8e",
   845 => x"1480f52d",
   846 => x"73708105",
   847 => x"5581b72d",
   848 => x"901480f5",
   849 => x"2d737081",
   850 => x"055581b7",
   851 => x"2d921480",
   852 => x"f52d7370",
   853 => x"81055581",
   854 => x"b72d9414",
   855 => x"80f52d73",
   856 => x"70810555",
   857 => x"81b72d96",
   858 => x"1480f52d",
   859 => x"73708105",
   860 => x"5581b72d",
   861 => x"981480f5",
   862 => x"2d737081",
   863 => x"055581b7",
   864 => x"2d9c1480",
   865 => x"f52d7370",
   866 => x"81055581",
   867 => x"b72d9e14",
   868 => x"80f52d73",
   869 => x"81b72d77",
   870 => x"bbbc0c80",
   871 => x"5372bc8c",
   872 => x"0c02a005",
   873 => x"0d0402cc",
   874 => x"050d7e60",
   875 => x"5e5a800b",
   876 => x"80c5f408",
   877 => x"80c5f808",
   878 => x"595c5680",
   879 => x"5880c5d4",
   880 => x"08782e81",
   881 => x"b038778f",
   882 => x"06a01757",
   883 => x"54738f38",
   884 => x"bfc45276",
   885 => x"51811757",
   886 => x"a5af2dbf",
   887 => x"c4568076",
   888 => x"80f52d56",
   889 => x"5474742e",
   890 => x"83388154",
   891 => x"7481e52e",
   892 => x"80f73881",
   893 => x"70750655",
   894 => x"5c73802e",
   895 => x"80eb388b",
   896 => x"1680f52d",
   897 => x"98065978",
   898 => x"80df388b",
   899 => x"537c5275",
   900 => x"5190d32d",
   901 => x"bc8c0880",
   902 => x"d0389c16",
   903 => x"0851a6cf",
   904 => x"2dbc8c08",
   905 => x"841b0c9a",
   906 => x"1680e02d",
   907 => x"51a6ff2d",
   908 => x"bc8c08bc",
   909 => x"8c08881c",
   910 => x"0cbc8c08",
   911 => x"555580c5",
   912 => x"d008802e",
   913 => x"98389416",
   914 => x"80e02d51",
   915 => x"a6ff2dbc",
   916 => x"8c08902b",
   917 => x"83fff00a",
   918 => x"06701651",
   919 => x"5473881b",
   920 => x"0c787a0c",
   921 => x"7b549dae",
   922 => x"04811858",
   923 => x"80c5d408",
   924 => x"7826fed2",
   925 => x"3880c5d0",
   926 => x"08802eb0",
   927 => x"387a5198",
   928 => x"802dbc8c",
   929 => x"08bc8c08",
   930 => x"80ffffff",
   931 => x"f806555b",
   932 => x"7380ffff",
   933 => x"fff82e94",
   934 => x"38bc8c08",
   935 => x"fe0580c5",
   936 => x"c8082980",
   937 => x"c5dc0805",
   938 => x"579bbb04",
   939 => x"805473bc",
   940 => x"8c0c02b4",
   941 => x"050d0402",
   942 => x"f4050d74",
   943 => x"70088105",
   944 => x"710c7008",
   945 => x"80c5cc08",
   946 => x"06535371",
   947 => x"8e388813",
   948 => x"08519880",
   949 => x"2dbc8c08",
   950 => x"88140c81",
   951 => x"0bbc8c0c",
   952 => x"028c050d",
   953 => x"0402f005",
   954 => x"0d758811",
   955 => x"08fe0580",
   956 => x"c5c80829",
   957 => x"80c5dc08",
   958 => x"11720880",
   959 => x"c5cc0806",
   960 => x"05795553",
   961 => x"5454a5af",
   962 => x"2d029005",
   963 => x"0d0402f0",
   964 => x"050d7588",
   965 => x"1108fe05",
   966 => x"80c5c808",
   967 => x"2980c5dc",
   968 => x"08117208",
   969 => x"80c5cc08",
   970 => x"06057955",
   971 => x"535454a3",
   972 => x"ef2d0290",
   973 => x"050d0402",
   974 => x"f4050dd4",
   975 => x"5281ff72",
   976 => x"0c710853",
   977 => x"81ff720c",
   978 => x"72882b83",
   979 => x"fe800672",
   980 => x"087081ff",
   981 => x"06515253",
   982 => x"81ff720c",
   983 => x"72710788",
   984 => x"2b720870",
   985 => x"81ff0651",
   986 => x"525381ff",
   987 => x"720c7271",
   988 => x"07882b72",
   989 => x"087081ff",
   990 => x"067207bc",
   991 => x"8c0c5253",
   992 => x"028c050d",
   993 => x"0402f405",
   994 => x"0d747671",
   995 => x"81ff06d4",
   996 => x"0c535380",
   997 => x"c6800885",
   998 => x"3871892b",
   999 => x"5271982a",
  1000 => x"d40c7190",
  1001 => x"2a7081ff",
  1002 => x"06d40c51",
  1003 => x"71882a70",
  1004 => x"81ff06d4",
  1005 => x"0c517181",
  1006 => x"ff06d40c",
  1007 => x"72902a70",
  1008 => x"81ff06d4",
  1009 => x"0c51d408",
  1010 => x"7081ff06",
  1011 => x"515182b8",
  1012 => x"bf527081",
  1013 => x"ff2e0981",
  1014 => x"06943881",
  1015 => x"ff0bd40c",
  1016 => x"d4087081",
  1017 => x"ff06ff14",
  1018 => x"54515171",
  1019 => x"e53870bc",
  1020 => x"8c0c028c",
  1021 => x"050d0402",
  1022 => x"fc050d81",
  1023 => x"c75181ff",
  1024 => x"0bd40cff",
  1025 => x"11517080",
  1026 => x"25f43802",
  1027 => x"84050d04",
  1028 => x"02f0050d",
  1029 => x"9ff72d8f",
  1030 => x"cf538052",
  1031 => x"87fc80f7",
  1032 => x"519f852d",
  1033 => x"bc8c0854",
  1034 => x"bc8c0881",
  1035 => x"2e098106",
  1036 => x"a33881ff",
  1037 => x"0bd40c82",
  1038 => x"0a52849c",
  1039 => x"80e9519f",
  1040 => x"852dbc8c",
  1041 => x"088b3881",
  1042 => x"ff0bd40c",
  1043 => x"7353a0da",
  1044 => x"049ff72d",
  1045 => x"ff135372",
  1046 => x"c13872bc",
  1047 => x"8c0c0290",
  1048 => x"050d0402",
  1049 => x"f4050d81",
  1050 => x"ff0bd40c",
  1051 => x"93538052",
  1052 => x"87fc80c1",
  1053 => x"519f852d",
  1054 => x"bc8c088b",
  1055 => x"3881ff0b",
  1056 => x"d40c8153",
  1057 => x"a190049f",
  1058 => x"f72dff13",
  1059 => x"5372df38",
  1060 => x"72bc8c0c",
  1061 => x"028c050d",
  1062 => x"0402f005",
  1063 => x"0d9ff72d",
  1064 => x"83aa5284",
  1065 => x"9c80c851",
  1066 => x"9f852dbc",
  1067 => x"8c08812e",
  1068 => x"09810692",
  1069 => x"389eb72d",
  1070 => x"bc8c0883",
  1071 => x"ffff0653",
  1072 => x"7283aa2e",
  1073 => x"9738a0e3",
  1074 => x"2da1d704",
  1075 => x"8154a2bc",
  1076 => x"04b8c451",
  1077 => x"85f22d80",
  1078 => x"54a2bc04",
  1079 => x"81ff0bd4",
  1080 => x"0cb153a0",
  1081 => x"902dbc8c",
  1082 => x"08802e80",
  1083 => x"c0388052",
  1084 => x"87fc80fa",
  1085 => x"519f852d",
  1086 => x"bc8c08b1",
  1087 => x"3881ff0b",
  1088 => x"d40cd408",
  1089 => x"5381ff0b",
  1090 => x"d40c81ff",
  1091 => x"0bd40c81",
  1092 => x"ff0bd40c",
  1093 => x"81ff0bd4",
  1094 => x"0c72862a",
  1095 => x"708106bc",
  1096 => x"8c085651",
  1097 => x"5372802e",
  1098 => x"9338a1cc",
  1099 => x"0472822e",
  1100 => x"ff9f38ff",
  1101 => x"135372ff",
  1102 => x"aa387254",
  1103 => x"73bc8c0c",
  1104 => x"0290050d",
  1105 => x"0402f005",
  1106 => x"0d810b80",
  1107 => x"c6800c84",
  1108 => x"54d00870",
  1109 => x"8f2a7081",
  1110 => x"06515153",
  1111 => x"72f33872",
  1112 => x"d00c9ff7",
  1113 => x"2db8d451",
  1114 => x"85f22dd0",
  1115 => x"08708f2a",
  1116 => x"70810651",
  1117 => x"515372f3",
  1118 => x"38810bd0",
  1119 => x"0cb15380",
  1120 => x"5284d480",
  1121 => x"c0519f85",
  1122 => x"2dbc8c08",
  1123 => x"812ea138",
  1124 => x"72822e09",
  1125 => x"81068c38",
  1126 => x"b8e05185",
  1127 => x"f22d8053",
  1128 => x"a3e604ff",
  1129 => x"135372d7",
  1130 => x"38ff1454",
  1131 => x"73ffa238",
  1132 => x"a1992dbc",
  1133 => x"8c0880c6",
  1134 => x"800cbc8c",
  1135 => x"088b3881",
  1136 => x"5287fc80",
  1137 => x"d0519f85",
  1138 => x"2d81ff0b",
  1139 => x"d40cd008",
  1140 => x"708f2a70",
  1141 => x"81065151",
  1142 => x"5372f338",
  1143 => x"72d00c81",
  1144 => x"ff0bd40c",
  1145 => x"815372bc",
  1146 => x"8c0c0290",
  1147 => x"050d0402",
  1148 => x"e8050d78",
  1149 => x"5681ff0b",
  1150 => x"d40cd008",
  1151 => x"708f2a70",
  1152 => x"81065151",
  1153 => x"5372f338",
  1154 => x"82810bd0",
  1155 => x"0c81ff0b",
  1156 => x"d40c7752",
  1157 => x"87fc80d8",
  1158 => x"519f852d",
  1159 => x"bc8c0880",
  1160 => x"2e8c38b8",
  1161 => x"f85185f2",
  1162 => x"2d8153a5",
  1163 => x"a60481ff",
  1164 => x"0bd40c81",
  1165 => x"fe0bd40c",
  1166 => x"80ff5575",
  1167 => x"70840557",
  1168 => x"0870982a",
  1169 => x"d40c7090",
  1170 => x"2c7081ff",
  1171 => x"06d40c54",
  1172 => x"70882c70",
  1173 => x"81ff06d4",
  1174 => x"0c547081",
  1175 => x"ff06d40c",
  1176 => x"54ff1555",
  1177 => x"748025d3",
  1178 => x"3881ff0b",
  1179 => x"d40c81ff",
  1180 => x"0bd40c81",
  1181 => x"ff0bd40c",
  1182 => x"868da054",
  1183 => x"81ff0bd4",
  1184 => x"0cd40881",
  1185 => x"ff065574",
  1186 => x"8738ff14",
  1187 => x"5473ed38",
  1188 => x"81ff0bd4",
  1189 => x"0cd00870",
  1190 => x"8f2a7081",
  1191 => x"06515153",
  1192 => x"72f33872",
  1193 => x"d00c72bc",
  1194 => x"8c0c0298",
  1195 => x"050d0402",
  1196 => x"e8050d78",
  1197 => x"55805681",
  1198 => x"ff0bd40c",
  1199 => x"d008708f",
  1200 => x"2a708106",
  1201 => x"51515372",
  1202 => x"f3388281",
  1203 => x"0bd00c81",
  1204 => x"ff0bd40c",
  1205 => x"775287fc",
  1206 => x"80d1519f",
  1207 => x"852d80db",
  1208 => x"c6df54bc",
  1209 => x"8c08802e",
  1210 => x"8a38b988",
  1211 => x"5185f22d",
  1212 => x"a6c60481",
  1213 => x"ff0bd40c",
  1214 => x"d4087081",
  1215 => x"ff065153",
  1216 => x"7281fe2e",
  1217 => x"0981069d",
  1218 => x"3880ff53",
  1219 => x"9eb72dbc",
  1220 => x"8c087570",
  1221 => x"8405570c",
  1222 => x"ff135372",
  1223 => x"8025ed38",
  1224 => x"8156a6ab",
  1225 => x"04ff1454",
  1226 => x"73c93881",
  1227 => x"ff0bd40c",
  1228 => x"81ff0bd4",
  1229 => x"0cd00870",
  1230 => x"8f2a7081",
  1231 => x"06515153",
  1232 => x"72f33872",
  1233 => x"d00c75bc",
  1234 => x"8c0c0298",
  1235 => x"050d0402",
  1236 => x"f4050d74",
  1237 => x"70882a83",
  1238 => x"fe800670",
  1239 => x"72982a07",
  1240 => x"72882b87",
  1241 => x"fc808006",
  1242 => x"73982b81",
  1243 => x"f00a0671",
  1244 => x"730707bc",
  1245 => x"8c0c5651",
  1246 => x"5351028c",
  1247 => x"050d0402",
  1248 => x"f8050d02",
  1249 => x"8e0580f5",
  1250 => x"2d74882b",
  1251 => x"077083ff",
  1252 => x"ff06bc8c",
  1253 => x"0c510288",
  1254 => x"050d0402",
  1255 => x"fc050d72",
  1256 => x"5180710c",
  1257 => x"800b8412",
  1258 => x"0c028405",
  1259 => x"0d0402f0",
  1260 => x"050d7570",
  1261 => x"08841208",
  1262 => x"535353ff",
  1263 => x"5471712e",
  1264 => x"a838aaf2",
  1265 => x"2d841308",
  1266 => x"70842914",
  1267 => x"88117008",
  1268 => x"7081ff06",
  1269 => x"84180881",
  1270 => x"11870684",
  1271 => x"1a0c5351",
  1272 => x"55515151",
  1273 => x"aaec2d71",
  1274 => x"5473bc8c",
  1275 => x"0c029005",
  1276 => x"0d0402f8",
  1277 => x"050daaf2",
  1278 => x"2de00870",
  1279 => x"8b2a7081",
  1280 => x"06515252",
  1281 => x"70802ea1",
  1282 => x"3880c684",
  1283 => x"08708429",
  1284 => x"80c68c05",
  1285 => x"7381ff06",
  1286 => x"710c5151",
  1287 => x"80c68408",
  1288 => x"81118706",
  1289 => x"80c6840c",
  1290 => x"51800b80",
  1291 => x"c6ac0caa",
  1292 => x"e52daaec",
  1293 => x"2d028805",
  1294 => x"0d0402fc",
  1295 => x"050daaf2",
  1296 => x"2d810b80",
  1297 => x"c6ac0caa",
  1298 => x"ec2d80c6",
  1299 => x"ac085170",
  1300 => x"f9380284",
  1301 => x"050d0402",
  1302 => x"fc050d80",
  1303 => x"c68451a7",
  1304 => x"9b2da7f2",
  1305 => x"51aae12d",
  1306 => x"aa8b2d02",
  1307 => x"84050d04",
  1308 => x"02f4050d",
  1309 => x"a9f204bc",
  1310 => x"8c0881f0",
  1311 => x"2e098106",
  1312 => x"8938810b",
  1313 => x"bc800ca9",
  1314 => x"f204bc8c",
  1315 => x"0881e02e",
  1316 => x"09810689",
  1317 => x"38810bbc",
  1318 => x"840ca9f2",
  1319 => x"04bc8c08",
  1320 => x"52bc8408",
  1321 => x"802e8838",
  1322 => x"bc8c0881",
  1323 => x"80055271",
  1324 => x"842c728f",
  1325 => x"065353bc",
  1326 => x"8008802e",
  1327 => x"99387284",
  1328 => x"29bbc005",
  1329 => x"72138171",
  1330 => x"2b700973",
  1331 => x"0806730c",
  1332 => x"515353a9",
  1333 => x"e8047284",
  1334 => x"29bbc005",
  1335 => x"72138371",
  1336 => x"2b720807",
  1337 => x"720c5353",
  1338 => x"800bbc84",
  1339 => x"0c800bbc",
  1340 => x"800c80c6",
  1341 => x"8451a7ae",
  1342 => x"2dbc8c08",
  1343 => x"ff24fef7",
  1344 => x"38800bbc",
  1345 => x"8c0c028c",
  1346 => x"050d0402",
  1347 => x"f8050dbb",
  1348 => x"c0528f51",
  1349 => x"80727084",
  1350 => x"05540cff",
  1351 => x"11517080",
  1352 => x"25f23802",
  1353 => x"88050d04",
  1354 => x"02f0050d",
  1355 => x"7551aaf2",
  1356 => x"2d70822c",
  1357 => x"fc06bbc0",
  1358 => x"1172109e",
  1359 => x"06710870",
  1360 => x"722a7083",
  1361 => x"0682742b",
  1362 => x"70097406",
  1363 => x"760c5451",
  1364 => x"56575351",
  1365 => x"53aaec2d",
  1366 => x"71bc8c0c",
  1367 => x"0290050d",
  1368 => x"0471980c",
  1369 => x"04ffb008",
  1370 => x"bc8c0c04",
  1371 => x"810bffb0",
  1372 => x"0c04800b",
  1373 => x"ffb00c04",
  1374 => x"02fc050d",
  1375 => x"810bbc88",
  1376 => x"0c815184",
  1377 => x"e62d0284",
  1378 => x"050d0402",
  1379 => x"fc050d80",
  1380 => x"0bbc880c",
  1381 => x"805184e6",
  1382 => x"2d028405",
  1383 => x"0d0402ec",
  1384 => x"050d7654",
  1385 => x"8052870b",
  1386 => x"881580f5",
  1387 => x"2d565374",
  1388 => x"72248338",
  1389 => x"a0537251",
  1390 => x"82ef2d81",
  1391 => x"128b1580",
  1392 => x"f52d5452",
  1393 => x"727225de",
  1394 => x"38029405",
  1395 => x"0d0402f0",
  1396 => x"050d80c6",
  1397 => x"bc085481",
  1398 => x"f82d800b",
  1399 => x"80c6c00c",
  1400 => x"7308802e",
  1401 => x"81843882",
  1402 => x"0bbca00c",
  1403 => x"80c6c008",
  1404 => x"8f06bc9c",
  1405 => x"0c730852",
  1406 => x"71832e96",
  1407 => x"38718326",
  1408 => x"89387181",
  1409 => x"2eaf38ac",
  1410 => x"d3047185",
  1411 => x"2e9f38ac",
  1412 => x"d3048814",
  1413 => x"80f52d84",
  1414 => x"1508b998",
  1415 => x"53545285",
  1416 => x"f22d7184",
  1417 => x"29137008",
  1418 => x"5252acd7",
  1419 => x"047351ab",
  1420 => x"9e2dacd3",
  1421 => x"0480c6b0",
  1422 => x"08881508",
  1423 => x"2c708106",
  1424 => x"51527180",
  1425 => x"2e8738b9",
  1426 => x"9c51acd0",
  1427 => x"04b9a051",
  1428 => x"85f22d84",
  1429 => x"14085185",
  1430 => x"f22d80c6",
  1431 => x"c0088105",
  1432 => x"80c6c00c",
  1433 => x"8c1454ab",
  1434 => x"e0040290",
  1435 => x"050d0471",
  1436 => x"80c6bc0c",
  1437 => x"abce2d80",
  1438 => x"c6c008ff",
  1439 => x"0580c6c4",
  1440 => x"0c0402e8",
  1441 => x"050d80c6",
  1442 => x"bc0880c6",
  1443 => x"c8085755",
  1444 => x"80f851aa",
  1445 => x"a82dbc8c",
  1446 => x"08812a70",
  1447 => x"81065152",
  1448 => x"719b3887",
  1449 => x"51aaa82d",
  1450 => x"bc8c0881",
  1451 => x"2a708106",
  1452 => x"51527180",
  1453 => x"2eb138ad",
  1454 => x"bd04a8f0",
  1455 => x"2d8751aa",
  1456 => x"a82dbc8c",
  1457 => x"08f438ad",
  1458 => x"cd04a8f0",
  1459 => x"2d80f851",
  1460 => x"aaa82dbc",
  1461 => x"8c08f338",
  1462 => x"bc880881",
  1463 => x"3270bc88",
  1464 => x"0c705252",
  1465 => x"84e62d80",
  1466 => x"0b80c6b4",
  1467 => x"0c800b80",
  1468 => x"c6b80cbc",
  1469 => x"880882fd",
  1470 => x"3880da51",
  1471 => x"aaa82dbc",
  1472 => x"8c08802e",
  1473 => x"8c3880c6",
  1474 => x"b4088180",
  1475 => x"0780c6b4",
  1476 => x"0c80d951",
  1477 => x"aaa82dbc",
  1478 => x"8c08802e",
  1479 => x"8c3880c6",
  1480 => x"b40880c0",
  1481 => x"0780c6b4",
  1482 => x"0c819451",
  1483 => x"aaa82dbc",
  1484 => x"8c08802e",
  1485 => x"8b3880c6",
  1486 => x"b4089007",
  1487 => x"80c6b40c",
  1488 => x"819151aa",
  1489 => x"a82dbc8c",
  1490 => x"08802e8b",
  1491 => x"3880c6b4",
  1492 => x"08a00780",
  1493 => x"c6b40c81",
  1494 => x"f551aaa8",
  1495 => x"2dbc8c08",
  1496 => x"802e8b38",
  1497 => x"80c6b408",
  1498 => x"810780c6",
  1499 => x"b40c81f2",
  1500 => x"51aaa82d",
  1501 => x"bc8c0880",
  1502 => x"2e8b3880",
  1503 => x"c6b40882",
  1504 => x"0780c6b4",
  1505 => x"0c81eb51",
  1506 => x"aaa82dbc",
  1507 => x"8c08802e",
  1508 => x"8b3880c6",
  1509 => x"b4088407",
  1510 => x"80c6b40c",
  1511 => x"81f451aa",
  1512 => x"a82dbc8c",
  1513 => x"08802e8b",
  1514 => x"3880c6b4",
  1515 => x"08880780",
  1516 => x"c6b40c80",
  1517 => x"d851aaa8",
  1518 => x"2dbc8c08",
  1519 => x"802e8c38",
  1520 => x"80c6b808",
  1521 => x"81800780",
  1522 => x"c6b80c92",
  1523 => x"51aaa82d",
  1524 => x"bc8c0880",
  1525 => x"2e8c3880",
  1526 => x"c6b80880",
  1527 => x"c00780c6",
  1528 => x"b80c9451",
  1529 => x"aaa82dbc",
  1530 => x"8c08802e",
  1531 => x"8b3880c6",
  1532 => x"b8089007",
  1533 => x"80c6b80c",
  1534 => x"9151aaa8",
  1535 => x"2dbc8c08",
  1536 => x"802e8b38",
  1537 => x"80c6b808",
  1538 => x"a00780c6",
  1539 => x"b80c9d51",
  1540 => x"aaa82dbc",
  1541 => x"8c08802e",
  1542 => x"8b3880c6",
  1543 => x"b8088107",
  1544 => x"80c6b80c",
  1545 => x"9b51aaa8",
  1546 => x"2dbc8c08",
  1547 => x"802e8b38",
  1548 => x"80c6b808",
  1549 => x"820780c6",
  1550 => x"b80c9c51",
  1551 => x"aaa82dbc",
  1552 => x"8c08802e",
  1553 => x"8b3880c6",
  1554 => x"b8088407",
  1555 => x"80c6b80c",
  1556 => x"a351aaa8",
  1557 => x"2dbc8c08",
  1558 => x"802e8b38",
  1559 => x"80c6b808",
  1560 => x"880780c6",
  1561 => x"b80c81fd",
  1562 => x"51aaa82d",
  1563 => x"81fa51aa",
  1564 => x"a82db6bd",
  1565 => x"0481f551",
  1566 => x"aaa82dbc",
  1567 => x"8c08812a",
  1568 => x"70810651",
  1569 => x"5271802e",
  1570 => x"b33880c6",
  1571 => x"c4085271",
  1572 => x"802e8a38",
  1573 => x"ff1280c6",
  1574 => x"c40cb1bc",
  1575 => x"0480c6c0",
  1576 => x"081080c6",
  1577 => x"c0080570",
  1578 => x"84291651",
  1579 => x"52881208",
  1580 => x"802e8938",
  1581 => x"ff518812",
  1582 => x"0852712d",
  1583 => x"81f251aa",
  1584 => x"a82dbc8c",
  1585 => x"08812a70",
  1586 => x"81065152",
  1587 => x"71802eb4",
  1588 => x"3880c6c0",
  1589 => x"08ff1180",
  1590 => x"c6c40856",
  1591 => x"53537372",
  1592 => x"258a3881",
  1593 => x"1480c6c4",
  1594 => x"0cb28404",
  1595 => x"72101370",
  1596 => x"84291651",
  1597 => x"52881208",
  1598 => x"802e8938",
  1599 => x"fe518812",
  1600 => x"0852712d",
  1601 => x"81fd51aa",
  1602 => x"a82dbc8c",
  1603 => x"08812a70",
  1604 => x"81065152",
  1605 => x"71802eb1",
  1606 => x"3880c6c4",
  1607 => x"08802e8a",
  1608 => x"38800b80",
  1609 => x"c6c40cb2",
  1610 => x"c90480c6",
  1611 => x"c0081080",
  1612 => x"c6c00805",
  1613 => x"70842916",
  1614 => x"51528812",
  1615 => x"08802e89",
  1616 => x"38fd5188",
  1617 => x"12085271",
  1618 => x"2d81fa51",
  1619 => x"aaa82dbc",
  1620 => x"8c08812a",
  1621 => x"70810651",
  1622 => x"5271802e",
  1623 => x"b13880c6",
  1624 => x"c008ff11",
  1625 => x"545280c6",
  1626 => x"c4087325",
  1627 => x"89387280",
  1628 => x"c6c40cb3",
  1629 => x"8e047110",
  1630 => x"12708429",
  1631 => x"16515288",
  1632 => x"1208802e",
  1633 => x"8938fc51",
  1634 => x"88120852",
  1635 => x"712d80c6",
  1636 => x"c4087053",
  1637 => x"5473802e",
  1638 => x"8a388c15",
  1639 => x"ff155555",
  1640 => x"b3950482",
  1641 => x"0bbca00c",
  1642 => x"718f06bc",
  1643 => x"9c0c81eb",
  1644 => x"51aaa82d",
  1645 => x"bc8c0881",
  1646 => x"2a708106",
  1647 => x"51527180",
  1648 => x"2ead3874",
  1649 => x"08852e09",
  1650 => x"8106a438",
  1651 => x"881580f5",
  1652 => x"2dff0552",
  1653 => x"71881681",
  1654 => x"b72d7198",
  1655 => x"2b527180",
  1656 => x"25883880",
  1657 => x"0b881681",
  1658 => x"b72d7451",
  1659 => x"ab9e2d81",
  1660 => x"f451aaa8",
  1661 => x"2dbc8c08",
  1662 => x"812a7081",
  1663 => x"06515271",
  1664 => x"802eb338",
  1665 => x"7408852e",
  1666 => x"098106aa",
  1667 => x"38881580",
  1668 => x"f52d8105",
  1669 => x"52718816",
  1670 => x"81b72d71",
  1671 => x"81ff068b",
  1672 => x"1680f52d",
  1673 => x"54527272",
  1674 => x"27873872",
  1675 => x"881681b7",
  1676 => x"2d7451ab",
  1677 => x"9e2d80da",
  1678 => x"51aaa82d",
  1679 => x"bc8c0881",
  1680 => x"2a708106",
  1681 => x"51527180",
  1682 => x"2e81ac38",
  1683 => x"80c6bc08",
  1684 => x"80c6c408",
  1685 => x"55537380",
  1686 => x"2e8a388c",
  1687 => x"13ff1555",
  1688 => x"53b4d604",
  1689 => x"72085271",
  1690 => x"822ea638",
  1691 => x"71822689",
  1692 => x"3871812e",
  1693 => x"aa38b5f7",
  1694 => x"0471832e",
  1695 => x"b4387184",
  1696 => x"2e098106",
  1697 => x"80f13888",
  1698 => x"130851ac",
  1699 => x"ef2db5f7",
  1700 => x"0480c6c4",
  1701 => x"08518813",
  1702 => x"0852712d",
  1703 => x"b5f70481",
  1704 => x"0b881408",
  1705 => x"2b80c6b0",
  1706 => x"083280c6",
  1707 => x"b00cb5cc",
  1708 => x"04881380",
  1709 => x"f52d8105",
  1710 => x"8b1480f5",
  1711 => x"2d535471",
  1712 => x"74248338",
  1713 => x"80547388",
  1714 => x"1481b72d",
  1715 => x"abce2db5",
  1716 => x"f7047508",
  1717 => x"802ea338",
  1718 => x"750851aa",
  1719 => x"a82dbc8c",
  1720 => x"08810652",
  1721 => x"71802e8c",
  1722 => x"3880c6c4",
  1723 => x"08518416",
  1724 => x"0852712d",
  1725 => x"88165675",
  1726 => x"d9388054",
  1727 => x"800bbca0",
  1728 => x"0c738f06",
  1729 => x"bc9c0ca0",
  1730 => x"527380c6",
  1731 => x"c4082e09",
  1732 => x"81069938",
  1733 => x"80c6c008",
  1734 => x"ff057432",
  1735 => x"70098105",
  1736 => x"7072079f",
  1737 => x"2a917131",
  1738 => x"51515353",
  1739 => x"715182ef",
  1740 => x"2d811454",
  1741 => x"8e7425c4",
  1742 => x"38bc8808",
  1743 => x"5271bc8c",
  1744 => x"0c029805",
  1745 => x"0d040000",
  1746 => x"00ffffff",
  1747 => x"ff00ffff",
  1748 => x"ffff00ff",
  1749 => x"ffffff00",
  1750 => x"52657365",
  1751 => x"74000000",
  1752 => x"53617665",
  1753 => x"20736574",
  1754 => x"74696e67",
  1755 => x"73000000",
  1756 => x"5363616e",
  1757 => x"6c696e65",
  1758 => x"73000000",
  1759 => x"4c6f6164",
  1760 => x"20524f4d",
  1761 => x"20100000",
  1762 => x"45786974",
  1763 => x"00000000",
  1764 => x"56474120",
  1765 => x"2d203331",
  1766 => x"4b487a2c",
  1767 => x"20363048",
  1768 => x"7a000000",
  1769 => x"5456202d",
  1770 => x"20343830",
  1771 => x"692c2036",
  1772 => x"30487a00",
  1773 => x"4261636b",
  1774 => x"00000000",
  1775 => x"46504741",
  1776 => x"47454e20",
  1777 => x"43464700",
  1778 => x"496e6974",
  1779 => x"69616c69",
  1780 => x"7a696e67",
  1781 => x"20534420",
  1782 => x"63617264",
  1783 => x"0a000000",
  1784 => x"424f4f54",
  1785 => x"20202020",
  1786 => x"47454e00",
  1787 => x"43617264",
  1788 => x"20696e69",
  1789 => x"74206661",
  1790 => x"696c6564",
  1791 => x"0a000000",
  1792 => x"4d425220",
  1793 => x"6661696c",
  1794 => x"0a000000",
  1795 => x"46415431",
  1796 => x"36202020",
  1797 => x"00000000",
  1798 => x"46415433",
  1799 => x"32202020",
  1800 => x"00000000",
  1801 => x"4e6f2070",
  1802 => x"61727469",
  1803 => x"74696f6e",
  1804 => x"20736967",
  1805 => x"0a000000",
  1806 => x"42616420",
  1807 => x"70617274",
  1808 => x"0a000000",
  1809 => x"53444843",
  1810 => x"20657272",
  1811 => x"6f72210a",
  1812 => x"00000000",
  1813 => x"53442069",
  1814 => x"6e69742e",
  1815 => x"2e2e0a00",
  1816 => x"53442063",
  1817 => x"61726420",
  1818 => x"72657365",
  1819 => x"74206661",
  1820 => x"696c6564",
  1821 => x"210a0000",
  1822 => x"57726974",
  1823 => x"65206661",
  1824 => x"696c6564",
  1825 => x"0a000000",
  1826 => x"52656164",
  1827 => x"20666169",
  1828 => x"6c65640a",
  1829 => x"00000000",
  1830 => x"16200000",
  1831 => x"14200000",
  1832 => x"15200000",
  1833 => x"00000002",
  1834 => x"00000002",
  1835 => x"00001b58",
  1836 => x"0000047f",
  1837 => x"00000002",
  1838 => x"00001b60",
  1839 => x"00000369",
  1840 => x"00000003",
  1841 => x"00001cfc",
  1842 => x"00000002",
  1843 => x"00000001",
  1844 => x"00001b70",
  1845 => x"00000001",
  1846 => x"00000002",
  1847 => x"00001b7c",
  1848 => x"00000719",
  1849 => x"00000002",
  1850 => x"00001b88",
  1851 => x"0000158b",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00001b90",
  1856 => x"00001ba4",
  1857 => x"00000002",
  1858 => x"00001e3c",
  1859 => x"0000050d",
  1860 => x"00000002",
  1861 => x"00001e5a",
  1862 => x"0000050d",
  1863 => x"00000002",
  1864 => x"00001e78",
  1865 => x"0000050d",
  1866 => x"00000002",
  1867 => x"00001e96",
  1868 => x"0000050d",
  1869 => x"00000002",
  1870 => x"00001eb4",
  1871 => x"0000050d",
  1872 => x"00000002",
  1873 => x"00001ed2",
  1874 => x"0000050d",
  1875 => x"00000002",
  1876 => x"00001ef0",
  1877 => x"0000050d",
  1878 => x"00000002",
  1879 => x"00001f0e",
  1880 => x"0000050d",
  1881 => x"00000002",
  1882 => x"00001f2c",
  1883 => x"0000050d",
  1884 => x"00000002",
  1885 => x"00001f4a",
  1886 => x"0000050d",
  1887 => x"00000002",
  1888 => x"00001f68",
  1889 => x"0000050d",
  1890 => x"00000002",
  1891 => x"00001f86",
  1892 => x"0000050d",
  1893 => x"00000002",
  1894 => x"00001fa4",
  1895 => x"0000050d",
  1896 => x"00000004",
  1897 => x"00001bb4",
  1898 => x"00001ca8",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"000006ad",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

