-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM1;

architecture arch of CtrlROM_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbe",
     9 => x"80080b0b",
    10 => x"0bbe8408",
    11 => x"0b0b0bbe",
    12 => x"88080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"be880c0b",
    16 => x"0b0bbe84",
    17 => x"0c0b0b0b",
    18 => x"be800c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb7c4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"be807080",
    57 => x"c8c0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518faf04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbe900c",
    65 => x"9f0bbe94",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"be9408ff",
    69 => x"05be940c",
    70 => x"be940880",
    71 => x"25eb38be",
    72 => x"9008ff05",
    73 => x"be900cbe",
    74 => x"90088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbe",
    94 => x"9008258f",
    95 => x"3882b32d",
    96 => x"be9008ff",
    97 => x"05be900c",
    98 => x"82f504be",
    99 => x"9008be94",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038be90",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"be940881",
   109 => x"05be940c",
   110 => x"be940851",
   111 => x"9f7125e2",
   112 => x"38800bbe",
   113 => x"940cbe90",
   114 => x"088105be",
   115 => x"900c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34be9408",
   120 => x"8105be94",
   121 => x"0cbe9408",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbe940c",
   125 => x"be900881",
   126 => x"05be900c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"be980cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbe",
   162 => x"980c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72be9808",
   167 => x"8407be98",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"bad00c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"be980852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c8a40cba",
   200 => x"f0718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"be800c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b8e852be",
   211 => x"9c519ca2",
   212 => x"2dbe8008",
   213 => x"802ea138",
   214 => x"80c1b852",
   215 => x"be9c519e",
   216 => x"e32d80c1",
   217 => x"b808bea8",
   218 => x"0c80c1b8",
   219 => x"08fec00c",
   220 => x"80c1b808",
   221 => x"5186932d",
   222 => x"0288050d",
   223 => x"0402f005",
   224 => x"0d805191",
   225 => x"f12db8e8",
   226 => x"52be9c51",
   227 => x"9ca22dbe",
   228 => x"8008802e",
   229 => x"a838bea8",
   230 => x"0880c1b8",
   231 => x"0c80c1bc",
   232 => x"5480fd53",
   233 => x"80747084",
   234 => x"05560cff",
   235 => x"13537280",
   236 => x"25f23880",
   237 => x"c1b852be",
   238 => x"9c519f8c",
   239 => x"2d029005",
   240 => x"0d0402d8",
   241 => x"050d800b",
   242 => x"bad40cbe",
   243 => x"a808fec0",
   244 => x"0c810bfe",
   245 => x"c40c840b",
   246 => x"fec40c7b",
   247 => x"52be9c51",
   248 => x"9ca22dbe",
   249 => x"800853be",
   250 => x"8008802e",
   251 => x"81b338be",
   252 => x"a0085580",
   253 => x"0bff1657",
   254 => x"5975792e",
   255 => x"8b388119",
   256 => x"76812a57",
   257 => x"5975f738",
   258 => x"f7195974",
   259 => x"b080802e",
   260 => x"09810689",
   261 => x"38820bfe",
   262 => x"dc0c88b4",
   263 => x"04749880",
   264 => x"802e0981",
   265 => x"06893881",
   266 => x"0bfedc0c",
   267 => x"88b40480",
   268 => x"0bfedc0c",
   269 => x"815a8075",
   270 => x"2580df38",
   271 => x"78527551",
   272 => x"84812d80",
   273 => x"c1b852be",
   274 => x"9c519ee3",
   275 => x"2dbe8008",
   276 => x"802ea838",
   277 => x"80c1b858",
   278 => x"83fc5777",
   279 => x"70840559",
   280 => x"087083ff",
   281 => x"ff067190",
   282 => x"2afec80c",
   283 => x"fec80cfc",
   284 => x"18585376",
   285 => x"8025e438",
   286 => x"898204be",
   287 => x"80085a84",
   288 => x"8055be9c",
   289 => x"519eb52d",
   290 => x"fc801581",
   291 => x"17575574",
   292 => x"8024ffa8",
   293 => x"3879802e",
   294 => x"8638820b",
   295 => x"bad40c79",
   296 => x"5372be80",
   297 => x"0c02a805",
   298 => x"0d0402fc",
   299 => x"050dac89",
   300 => x"2dfec451",
   301 => x"81710c82",
   302 => x"710c0284",
   303 => x"050d0402",
   304 => x"f4050d74",
   305 => x"76785354",
   306 => x"52807125",
   307 => x"97387270",
   308 => x"81055480",
   309 => x"f52d7270",
   310 => x"81055481",
   311 => x"b72dff11",
   312 => x"5170eb38",
   313 => x"807281b7",
   314 => x"2d028c05",
   315 => x"0d0402e8",
   316 => x"050d7756",
   317 => x"80705654",
   318 => x"737624b3",
   319 => x"3880c7c8",
   320 => x"08742eab",
   321 => x"38735199",
   322 => x"eb2dbe80",
   323 => x"08be8008",
   324 => x"09810570",
   325 => x"be800807",
   326 => x"9f2a7705",
   327 => x"81175757",
   328 => x"53537476",
   329 => x"24893880",
   330 => x"c7c80874",
   331 => x"26d73872",
   332 => x"be800c02",
   333 => x"98050d04",
   334 => x"02f4050d",
   335 => x"bcfc0815",
   336 => x"5189ee2d",
   337 => x"be800880",
   338 => x"2eaa388b",
   339 => x"53be8008",
   340 => x"5280c5b8",
   341 => x"5189bf2d",
   342 => x"80c5b851",
   343 => x"87c22dbe",
   344 => x"8008802e",
   345 => x"8f38bad8",
   346 => x"51aded2d",
   347 => x"ac892d80",
   348 => x"518aff04",
   349 => x"bd8051ad",
   350 => x"ed2dabf6",
   351 => x"2d815184",
   352 => x"e62d028c",
   353 => x"050d0402",
   354 => x"dc050d80",
   355 => x"705a5574",
   356 => x"bcfc0825",
   357 => x"b13880c7",
   358 => x"c808752e",
   359 => x"a9387851",
   360 => x"99eb2dbe",
   361 => x"80080981",
   362 => x"0570be80",
   363 => x"08079f2a",
   364 => x"7605811b",
   365 => x"5b565474",
   366 => x"bcfc0825",
   367 => x"893880c7",
   368 => x"c8087926",
   369 => x"d9388055",
   370 => x"7880c7c8",
   371 => x"082781d0",
   372 => x"38785199",
   373 => x"eb2dbe80",
   374 => x"08802e81",
   375 => x"a538be80",
   376 => x"088b0580",
   377 => x"f52d7084",
   378 => x"2a708106",
   379 => x"77107884",
   380 => x"2b80c5b8",
   381 => x"0b80f52d",
   382 => x"5c5c5351",
   383 => x"55567380",
   384 => x"2e80c738",
   385 => x"7416822b",
   386 => x"8dc30bbb",
   387 => x"d0120c54",
   388 => x"77753110",
   389 => x"beb01155",
   390 => x"56907470",
   391 => x"81055681",
   392 => x"b72da074",
   393 => x"81b72d76",
   394 => x"81ff0681",
   395 => x"16585473",
   396 => x"802e8a38",
   397 => x"9c5380c5",
   398 => x"b8528cc3",
   399 => x"048b53be",
   400 => x"800852be",
   401 => x"b216518c",
   402 => x"fa047416",
   403 => x"822b8ab8",
   404 => x"0bbbd012",
   405 => x"0c547681",
   406 => x"ff068116",
   407 => x"58547380",
   408 => x"2e8a389c",
   409 => x"5380c5b8",
   410 => x"528cf204",
   411 => x"8b53be80",
   412 => x"08527775",
   413 => x"3110beb0",
   414 => x"05517655",
   415 => x"89bf2d8d",
   416 => x"95047490",
   417 => x"29753170",
   418 => x"10beb005",
   419 => x"5154be80",
   420 => x"087481b7",
   421 => x"2d811959",
   422 => x"748b24a2",
   423 => x"388bc804",
   424 => x"74902975",
   425 => x"317010be",
   426 => x"b0058c77",
   427 => x"31575154",
   428 => x"807481b7",
   429 => x"2d9e14ff",
   430 => x"16565474",
   431 => x"f33802a4",
   432 => x"050d0402",
   433 => x"fc050dbc",
   434 => x"fc081351",
   435 => x"89ee2dbe",
   436 => x"8008802e",
   437 => x"8838be80",
   438 => x"085191f1",
   439 => x"2d800bbc",
   440 => x"fc0c8b87",
   441 => x"2daccc2d",
   442 => x"0284050d",
   443 => x"0402fc05",
   444 => x"0d725170",
   445 => x"fd2ead38",
   446 => x"70fd248a",
   447 => x"3870fc2e",
   448 => x"80c4388e",
   449 => x"ce0470fe",
   450 => x"2eb13870",
   451 => x"ff2e0981",
   452 => x"06bc38bc",
   453 => x"fc085170",
   454 => x"802eb338",
   455 => x"ff11bcfc",
   456 => x"0c8ece04",
   457 => x"bcfc08f0",
   458 => x"0570bcfc",
   459 => x"0c517080",
   460 => x"259c3880",
   461 => x"0bbcfc0c",
   462 => x"8ece04bc",
   463 => x"fc088105",
   464 => x"bcfc0c8e",
   465 => x"ce04bcfc",
   466 => x"089005bc",
   467 => x"fc0c8b87",
   468 => x"2daccc2d",
   469 => x"0284050d",
   470 => x"0402fc05",
   471 => x"0d800bbc",
   472 => x"fc0c8b87",
   473 => x"2dbbc851",
   474 => x"aded2d02",
   475 => x"84050d04",
   476 => x"02f8050d",
   477 => x"80c8a408",
   478 => x"8206baf8",
   479 => x"0b80f52d",
   480 => x"52527080",
   481 => x"2e853871",
   482 => x"810752bb",
   483 => x"900b80f5",
   484 => x"2d517080",
   485 => x"2e853871",
   486 => x"840752be",
   487 => x"ac08802e",
   488 => x"85387190",
   489 => x"075271be",
   490 => x"800c0288",
   491 => x"050d0402",
   492 => x"f4050d81",
   493 => x"0bbeac0c",
   494 => x"800bbad4",
   495 => x"0c905186",
   496 => x"932d810b",
   497 => x"fec40c84",
   498 => x"0bfec40c",
   499 => x"830bfecc",
   500 => x"0cb8f451",
   501 => x"85f22d84",
   502 => x"52a3c32d",
   503 => x"93922dbe",
   504 => x"8008802e",
   505 => x"8638fe52",
   506 => x"8ff304ff",
   507 => x"12527180",
   508 => x"24e73871",
   509 => x"802e81ab",
   510 => x"38a9d52d",
   511 => x"abea2da9",
   512 => x"b82da9b8",
   513 => x"2d81f82d",
   514 => x"815184e6",
   515 => x"2da9b82d",
   516 => x"a9b82d81",
   517 => x"5184e62d",
   518 => x"86c42db9",
   519 => x"8c5187c2",
   520 => x"2dbe8008",
   521 => x"802e9438",
   522 => x"bad851ad",
   523 => x"ed2d8051",
   524 => x"84e62d82",
   525 => x"0bbad40c",
   526 => x"90c504be",
   527 => x"8008518e",
   528 => x"d92dabf6",
   529 => x"2da9ee2d",
   530 => x"ae802dbe",
   531 => x"800880c8",
   532 => x"a808882b",
   533 => x"80c8ac08",
   534 => x"07fed80c",
   535 => x"538ef02d",
   536 => x"be8008be",
   537 => x"a8082ea2",
   538 => x"38be8008",
   539 => x"bea80cbe",
   540 => x"8008fec0",
   541 => x"0c845272",
   542 => x"5184e62d",
   543 => x"a9b82da9",
   544 => x"b82dff12",
   545 => x"52718025",
   546 => x"ee387280",
   547 => x"2e8c38ba",
   548 => x"d4088807",
   549 => x"fec40c90",
   550 => x"c504bad4",
   551 => x"08fec40c",
   552 => x"90c504b9",
   553 => x"985185f2",
   554 => x"2d800bbe",
   555 => x"800c028c",
   556 => x"050d0402",
   557 => x"e8050d77",
   558 => x"797b5855",
   559 => x"55805372",
   560 => x"7625a338",
   561 => x"74708105",
   562 => x"5680f52d",
   563 => x"74708105",
   564 => x"5680f52d",
   565 => x"52527171",
   566 => x"2e863881",
   567 => x"5191e804",
   568 => x"81135391",
   569 => x"bf048051",
   570 => x"70be800c",
   571 => x"0298050d",
   572 => x"0402ec05",
   573 => x"0d765574",
   574 => x"802ebe38",
   575 => x"9a1580e0",
   576 => x"2d51a7fd",
   577 => x"2dbe8008",
   578 => x"be800880",
   579 => x"c7e80cbe",
   580 => x"80085454",
   581 => x"80c7c408",
   582 => x"802e9938",
   583 => x"941580e0",
   584 => x"2d51a7fd",
   585 => x"2dbe8008",
   586 => x"902b83ff",
   587 => x"f00a0670",
   588 => x"75075153",
   589 => x"7280c7e8",
   590 => x"0c80c7e8",
   591 => x"08537280",
   592 => x"2e9d3880",
   593 => x"c7bc08fe",
   594 => x"14712980",
   595 => x"c7d00805",
   596 => x"80c7ec0c",
   597 => x"70842b80",
   598 => x"c7c80c54",
   599 => x"938d0480",
   600 => x"c7d40880",
   601 => x"c7e80c80",
   602 => x"c7d80880",
   603 => x"c7ec0c80",
   604 => x"c7c40880",
   605 => x"2e8b3880",
   606 => x"c7bc0884",
   607 => x"2b539388",
   608 => x"0480c7dc",
   609 => x"08842b53",
   610 => x"7280c7c8",
   611 => x"0c029405",
   612 => x"0d0402d8",
   613 => x"050d800b",
   614 => x"80c7c40c",
   615 => x"80c1b852",
   616 => x"8051a6ad",
   617 => x"2dbe8008",
   618 => x"54be8008",
   619 => x"8c38b9ac",
   620 => x"5185f22d",
   621 => x"735598ee",
   622 => x"04805681",
   623 => x"0b80c7f0",
   624 => x"0c8853b9",
   625 => x"b85280c1",
   626 => x"ee5191b3",
   627 => x"2dbe8008",
   628 => x"762e0981",
   629 => x"068838be",
   630 => x"800880c7",
   631 => x"f00c8853",
   632 => x"b9c45280",
   633 => x"c28a5191",
   634 => x"b32dbe80",
   635 => x"088838be",
   636 => x"800880c7",
   637 => x"f00c80c7",
   638 => x"f008802e",
   639 => x"80fd3880",
   640 => x"c4fe0b80",
   641 => x"f52d80c4",
   642 => x"ff0b80f5",
   643 => x"2d71982b",
   644 => x"71902b07",
   645 => x"80c5800b",
   646 => x"80f52d70",
   647 => x"882b7207",
   648 => x"80c5810b",
   649 => x"80f52d71",
   650 => x"0780c5b6",
   651 => x"0b80f52d",
   652 => x"80c5b70b",
   653 => x"80f52d71",
   654 => x"882b0753",
   655 => x"5f54525a",
   656 => x"56575573",
   657 => x"81abaa2e",
   658 => x"0981068d",
   659 => x"387551a7",
   660 => x"cd2dbe80",
   661 => x"085694e6",
   662 => x"047382d4",
   663 => x"d52e8738",
   664 => x"b9d05195",
   665 => x"ab0480c1",
   666 => x"b8527551",
   667 => x"a6ad2dbe",
   668 => x"800855be",
   669 => x"8008802e",
   670 => x"83f43888",
   671 => x"53b9c452",
   672 => x"80c28a51",
   673 => x"91b32dbe",
   674 => x"80088a38",
   675 => x"810b80c7",
   676 => x"c40c95b1",
   677 => x"048853b9",
   678 => x"b85280c1",
   679 => x"ee5191b3",
   680 => x"2dbe8008",
   681 => x"802e8a38",
   682 => x"b9e45185",
   683 => x"f22d9690",
   684 => x"0480c5b6",
   685 => x"0b80f52d",
   686 => x"547380d5",
   687 => x"2e098106",
   688 => x"80ce3880",
   689 => x"c5b70b80",
   690 => x"f52d5473",
   691 => x"81aa2e09",
   692 => x"8106bd38",
   693 => x"800b80c1",
   694 => x"b80b80f5",
   695 => x"2d565474",
   696 => x"81e92e83",
   697 => x"38815474",
   698 => x"81eb2e8c",
   699 => x"38805573",
   700 => x"752e0981",
   701 => x"0682f738",
   702 => x"80c1c30b",
   703 => x"80f52d55",
   704 => x"748e3880",
   705 => x"c1c40b80",
   706 => x"f52d5473",
   707 => x"822e8638",
   708 => x"805598ee",
   709 => x"0480c1c5",
   710 => x"0b80f52d",
   711 => x"7080c7bc",
   712 => x"0cff0580",
   713 => x"c7c00c80",
   714 => x"c1c60b80",
   715 => x"f52d80c1",
   716 => x"c70b80f5",
   717 => x"2d587605",
   718 => x"77828029",
   719 => x"057080c7",
   720 => x"cc0c80c1",
   721 => x"c80b80f5",
   722 => x"2d7080c7",
   723 => x"e00c80c7",
   724 => x"c4085957",
   725 => x"5876802e",
   726 => x"81b53888",
   727 => x"53b9c452",
   728 => x"80c28a51",
   729 => x"91b32dbe",
   730 => x"80088282",
   731 => x"3880c7bc",
   732 => x"0870842b",
   733 => x"80c7c80c",
   734 => x"7080c7dc",
   735 => x"0c80c1dd",
   736 => x"0b80f52d",
   737 => x"80c1dc0b",
   738 => x"80f52d71",
   739 => x"82802905",
   740 => x"80c1de0b",
   741 => x"80f52d70",
   742 => x"84808029",
   743 => x"1280c1df",
   744 => x"0b80f52d",
   745 => x"7081800a",
   746 => x"29127080",
   747 => x"c7e40c80",
   748 => x"c7e00871",
   749 => x"2980c7cc",
   750 => x"08057080",
   751 => x"c7d00c80",
   752 => x"c1e50b80",
   753 => x"f52d80c1",
   754 => x"e40b80f5",
   755 => x"2d718280",
   756 => x"290580c1",
   757 => x"e60b80f5",
   758 => x"2d708480",
   759 => x"80291280",
   760 => x"c1e70b80",
   761 => x"f52d7098",
   762 => x"2b81f00a",
   763 => x"06720570",
   764 => x"80c7d40c",
   765 => x"fe117e29",
   766 => x"770580c7",
   767 => x"d80c5259",
   768 => x"5243545e",
   769 => x"51525952",
   770 => x"5d575957",
   771 => x"98e70480",
   772 => x"c1ca0b80",
   773 => x"f52d80c1",
   774 => x"c90b80f5",
   775 => x"2d718280",
   776 => x"29057080",
   777 => x"c7c80c70",
   778 => x"a02983ff",
   779 => x"0570892a",
   780 => x"7080c7dc",
   781 => x"0c80c1cf",
   782 => x"0b80f52d",
   783 => x"80c1ce0b",
   784 => x"80f52d71",
   785 => x"82802905",
   786 => x"7080c7e4",
   787 => x"0c7b7129",
   788 => x"1e7080c7",
   789 => x"d80c7d80",
   790 => x"c7d40c73",
   791 => x"0580c7d0",
   792 => x"0c555e51",
   793 => x"51555580",
   794 => x"5191f12d",
   795 => x"815574be",
   796 => x"800c02a8",
   797 => x"050d0402",
   798 => x"ec050d76",
   799 => x"70872c71",
   800 => x"80ff0655",
   801 => x"565480c7",
   802 => x"c4088a38",
   803 => x"73882c74",
   804 => x"81ff0654",
   805 => x"5580c1b8",
   806 => x"5280c7cc",
   807 => x"081551a6",
   808 => x"ad2dbe80",
   809 => x"0854be80",
   810 => x"08802eb6",
   811 => x"3880c7c4",
   812 => x"08802e99",
   813 => x"38728429",
   814 => x"80c1b805",
   815 => x"70085253",
   816 => x"a7cd2dbe",
   817 => x"8008f00a",
   818 => x"065399e0",
   819 => x"04721080",
   820 => x"c1b80570",
   821 => x"80e02d52",
   822 => x"53a7fd2d",
   823 => x"be800853",
   824 => x"725473be",
   825 => x"800c0294",
   826 => x"050d0402",
   827 => x"e0050d79",
   828 => x"70842c80",
   829 => x"c7ec0805",
   830 => x"718f0652",
   831 => x"5553728a",
   832 => x"3880c1b8",
   833 => x"527351a6",
   834 => x"ad2d72a0",
   835 => x"2980c1b8",
   836 => x"05548074",
   837 => x"80f52d56",
   838 => x"5374732e",
   839 => x"83388153",
   840 => x"7481e52e",
   841 => x"81f13881",
   842 => x"70740654",
   843 => x"5872802e",
   844 => x"81e5388b",
   845 => x"1480f52d",
   846 => x"70832a79",
   847 => x"06585676",
   848 => x"9938bdb0",
   849 => x"08537289",
   850 => x"387280c5",
   851 => x"b80b81b7",
   852 => x"2d76bdb0",
   853 => x"0c73539c",
   854 => x"9904758f",
   855 => x"2e098106",
   856 => x"81b53874",
   857 => x"9f068d29",
   858 => x"80c5ab11",
   859 => x"51538114",
   860 => x"80f52d73",
   861 => x"70810555",
   862 => x"81b72d83",
   863 => x"1480f52d",
   864 => x"73708105",
   865 => x"5581b72d",
   866 => x"851480f5",
   867 => x"2d737081",
   868 => x"055581b7",
   869 => x"2d871480",
   870 => x"f52d7370",
   871 => x"81055581",
   872 => x"b72d8914",
   873 => x"80f52d73",
   874 => x"70810555",
   875 => x"81b72d8e",
   876 => x"1480f52d",
   877 => x"73708105",
   878 => x"5581b72d",
   879 => x"901480f5",
   880 => x"2d737081",
   881 => x"055581b7",
   882 => x"2d921480",
   883 => x"f52d7370",
   884 => x"81055581",
   885 => x"b72d9414",
   886 => x"80f52d73",
   887 => x"70810555",
   888 => x"81b72d96",
   889 => x"1480f52d",
   890 => x"73708105",
   891 => x"5581b72d",
   892 => x"981480f5",
   893 => x"2d737081",
   894 => x"055581b7",
   895 => x"2d9c1480",
   896 => x"f52d7370",
   897 => x"81055581",
   898 => x"b72d9e14",
   899 => x"80f52d73",
   900 => x"81b72d77",
   901 => x"bdb00c80",
   902 => x"5372be80",
   903 => x"0c02a005",
   904 => x"0d0402cc",
   905 => x"050d7e60",
   906 => x"5e5a800b",
   907 => x"80c7e808",
   908 => x"80c7ec08",
   909 => x"595c5680",
   910 => x"5880c7c8",
   911 => x"08782e81",
   912 => x"b238778f",
   913 => x"06a01757",
   914 => x"54739138",
   915 => x"80c1b852",
   916 => x"76518117",
   917 => x"57a6ad2d",
   918 => x"80c1b856",
   919 => x"807680f5",
   920 => x"2d565474",
   921 => x"742e8338",
   922 => x"81547481",
   923 => x"e52e80f7",
   924 => x"38817075",
   925 => x"06555c73",
   926 => x"802e80eb",
   927 => x"388b1680",
   928 => x"f52d9806",
   929 => x"597880df",
   930 => x"388b537c",
   931 => x"52755191",
   932 => x"b32dbe80",
   933 => x"0880d038",
   934 => x"9c160851",
   935 => x"a7cd2dbe",
   936 => x"8008841b",
   937 => x"0c9a1680",
   938 => x"e02d51a7",
   939 => x"fd2dbe80",
   940 => x"08be8008",
   941 => x"881c0cbe",
   942 => x"80085555",
   943 => x"80c7c408",
   944 => x"802e9838",
   945 => x"941680e0",
   946 => x"2d51a7fd",
   947 => x"2dbe8008",
   948 => x"902b83ff",
   949 => x"f00a0670",
   950 => x"16515473",
   951 => x"881b0c78",
   952 => x"7a0c7b54",
   953 => x"9eac0481",
   954 => x"185880c7",
   955 => x"c8087826",
   956 => x"fed03880",
   957 => x"c7c40880",
   958 => x"2eb0387a",
   959 => x"5198f72d",
   960 => x"be8008be",
   961 => x"800880ff",
   962 => x"fffff806",
   963 => x"555b7380",
   964 => x"fffffff8",
   965 => x"2e9438be",
   966 => x"8008fe05",
   967 => x"80c7bc08",
   968 => x"2980c7d0",
   969 => x"0805579c",
   970 => x"b7048054",
   971 => x"73be800c",
   972 => x"02b4050d",
   973 => x"0402f405",
   974 => x"0d747008",
   975 => x"8105710c",
   976 => x"700880c7",
   977 => x"c0080653",
   978 => x"53718e38",
   979 => x"88130851",
   980 => x"98f72dbe",
   981 => x"80088814",
   982 => x"0c810bbe",
   983 => x"800c028c",
   984 => x"050d0402",
   985 => x"f0050d75",
   986 => x"881108fe",
   987 => x"0580c7bc",
   988 => x"082980c7",
   989 => x"d0081172",
   990 => x"0880c7c0",
   991 => x"08060579",
   992 => x"55535454",
   993 => x"a6ad2d02",
   994 => x"90050d04",
   995 => x"02f0050d",
   996 => x"75881108",
   997 => x"fe0580c7",
   998 => x"bc082980",
   999 => x"c7d00811",
  1000 => x"720880c7",
  1001 => x"c0080605",
  1002 => x"79555354",
  1003 => x"54a4ed2d",
  1004 => x"0290050d",
  1005 => x"0402f405",
  1006 => x"0dd45281",
  1007 => x"ff720c71",
  1008 => x"085381ff",
  1009 => x"720c7288",
  1010 => x"2b83fe80",
  1011 => x"06720870",
  1012 => x"81ff0651",
  1013 => x"525381ff",
  1014 => x"720c7271",
  1015 => x"07882b72",
  1016 => x"087081ff",
  1017 => x"06515253",
  1018 => x"81ff720c",
  1019 => x"72710788",
  1020 => x"2b720870",
  1021 => x"81ff0672",
  1022 => x"07be800c",
  1023 => x"5253028c",
  1024 => x"050d0402",
  1025 => x"f4050d74",
  1026 => x"767181ff",
  1027 => x"06d40c53",
  1028 => x"5380c7f4",
  1029 => x"08853871",
  1030 => x"892b5271",
  1031 => x"982ad40c",
  1032 => x"71902a70",
  1033 => x"81ff06d4",
  1034 => x"0c517188",
  1035 => x"2a7081ff",
  1036 => x"06d40c51",
  1037 => x"7181ff06",
  1038 => x"d40c7290",
  1039 => x"2a7081ff",
  1040 => x"06d40c51",
  1041 => x"d4087081",
  1042 => x"ff065151",
  1043 => x"82b8bf52",
  1044 => x"7081ff2e",
  1045 => x"09810694",
  1046 => x"3881ff0b",
  1047 => x"d40cd408",
  1048 => x"7081ff06",
  1049 => x"ff145451",
  1050 => x"5171e538",
  1051 => x"70be800c",
  1052 => x"028c050d",
  1053 => x"0402fc05",
  1054 => x"0d81c751",
  1055 => x"81ff0bd4",
  1056 => x"0cff1151",
  1057 => x"708025f4",
  1058 => x"38028405",
  1059 => x"0d0402f0",
  1060 => x"050da0f5",
  1061 => x"2d8fcf53",
  1062 => x"805287fc",
  1063 => x"80f751a0",
  1064 => x"832dbe80",
  1065 => x"0854be80",
  1066 => x"08812e09",
  1067 => x"8106a338",
  1068 => x"81ff0bd4",
  1069 => x"0c820a52",
  1070 => x"849c80e9",
  1071 => x"51a0832d",
  1072 => x"be80088b",
  1073 => x"3881ff0b",
  1074 => x"d40c7353",
  1075 => x"a1d804a0",
  1076 => x"f52dff13",
  1077 => x"5372c138",
  1078 => x"72be800c",
  1079 => x"0290050d",
  1080 => x"0402f405",
  1081 => x"0d81ff0b",
  1082 => x"d40c9353",
  1083 => x"805287fc",
  1084 => x"80c151a0",
  1085 => x"832dbe80",
  1086 => x"088b3881",
  1087 => x"ff0bd40c",
  1088 => x"8153a28e",
  1089 => x"04a0f52d",
  1090 => x"ff135372",
  1091 => x"df3872be",
  1092 => x"800c028c",
  1093 => x"050d0402",
  1094 => x"f0050da0",
  1095 => x"f52d83aa",
  1096 => x"52849c80",
  1097 => x"c851a083",
  1098 => x"2dbe8008",
  1099 => x"812e0981",
  1100 => x"0692389f",
  1101 => x"b52dbe80",
  1102 => x"0883ffff",
  1103 => x"06537283",
  1104 => x"aa2e9738",
  1105 => x"a1e12da2",
  1106 => x"d5048154",
  1107 => x"a3ba04b9",
  1108 => x"f05185f2",
  1109 => x"2d8054a3",
  1110 => x"ba0481ff",
  1111 => x"0bd40cb1",
  1112 => x"53a18e2d",
  1113 => x"be800880",
  1114 => x"2e80c038",
  1115 => x"805287fc",
  1116 => x"80fa51a0",
  1117 => x"832dbe80",
  1118 => x"08b13881",
  1119 => x"ff0bd40c",
  1120 => x"d4085381",
  1121 => x"ff0bd40c",
  1122 => x"81ff0bd4",
  1123 => x"0c81ff0b",
  1124 => x"d40c81ff",
  1125 => x"0bd40c72",
  1126 => x"862a7081",
  1127 => x"06be8008",
  1128 => x"56515372",
  1129 => x"802e9338",
  1130 => x"a2ca0472",
  1131 => x"822eff9f",
  1132 => x"38ff1353",
  1133 => x"72ffaa38",
  1134 => x"725473be",
  1135 => x"800c0290",
  1136 => x"050d0402",
  1137 => x"f0050d81",
  1138 => x"0b80c7f4",
  1139 => x"0c8454d0",
  1140 => x"08708f2a",
  1141 => x"70810651",
  1142 => x"515372f3",
  1143 => x"3872d00c",
  1144 => x"a0f52dba",
  1145 => x"805185f2",
  1146 => x"2dd00870",
  1147 => x"8f2a7081",
  1148 => x"06515153",
  1149 => x"72f33881",
  1150 => x"0bd00cb1",
  1151 => x"53805284",
  1152 => x"d480c051",
  1153 => x"a0832dbe",
  1154 => x"8008812e",
  1155 => x"a1387282",
  1156 => x"2e098106",
  1157 => x"8c38ba8c",
  1158 => x"5185f22d",
  1159 => x"8053a4e4",
  1160 => x"04ff1353",
  1161 => x"72d738ff",
  1162 => x"145473ff",
  1163 => x"a238a297",
  1164 => x"2dbe8008",
  1165 => x"80c7f40c",
  1166 => x"be80088b",
  1167 => x"38815287",
  1168 => x"fc80d051",
  1169 => x"a0832d81",
  1170 => x"ff0bd40c",
  1171 => x"d008708f",
  1172 => x"2a708106",
  1173 => x"51515372",
  1174 => x"f33872d0",
  1175 => x"0c81ff0b",
  1176 => x"d40c8153",
  1177 => x"72be800c",
  1178 => x"0290050d",
  1179 => x"0402e805",
  1180 => x"0d785681",
  1181 => x"ff0bd40c",
  1182 => x"d008708f",
  1183 => x"2a708106",
  1184 => x"51515372",
  1185 => x"f3388281",
  1186 => x"0bd00c81",
  1187 => x"ff0bd40c",
  1188 => x"775287fc",
  1189 => x"80d851a0",
  1190 => x"832dbe80",
  1191 => x"08802e8c",
  1192 => x"38baa451",
  1193 => x"85f22d81",
  1194 => x"53a6a404",
  1195 => x"81ff0bd4",
  1196 => x"0c81fe0b",
  1197 => x"d40c80ff",
  1198 => x"55757084",
  1199 => x"05570870",
  1200 => x"982ad40c",
  1201 => x"70902c70",
  1202 => x"81ff06d4",
  1203 => x"0c547088",
  1204 => x"2c7081ff",
  1205 => x"06d40c54",
  1206 => x"7081ff06",
  1207 => x"d40c54ff",
  1208 => x"15557480",
  1209 => x"25d33881",
  1210 => x"ff0bd40c",
  1211 => x"81ff0bd4",
  1212 => x"0c81ff0b",
  1213 => x"d40c868d",
  1214 => x"a05481ff",
  1215 => x"0bd40cd4",
  1216 => x"0881ff06",
  1217 => x"55748738",
  1218 => x"ff145473",
  1219 => x"ed3881ff",
  1220 => x"0bd40cd0",
  1221 => x"08708f2a",
  1222 => x"70810651",
  1223 => x"515372f3",
  1224 => x"3872d00c",
  1225 => x"72be800c",
  1226 => x"0298050d",
  1227 => x"0402e805",
  1228 => x"0d785580",
  1229 => x"5681ff0b",
  1230 => x"d40cd008",
  1231 => x"708f2a70",
  1232 => x"81065151",
  1233 => x"5372f338",
  1234 => x"82810bd0",
  1235 => x"0c81ff0b",
  1236 => x"d40c7752",
  1237 => x"87fc80d1",
  1238 => x"51a0832d",
  1239 => x"80dbc6df",
  1240 => x"54be8008",
  1241 => x"802e8a38",
  1242 => x"bab45185",
  1243 => x"f22da7c4",
  1244 => x"0481ff0b",
  1245 => x"d40cd408",
  1246 => x"7081ff06",
  1247 => x"51537281",
  1248 => x"fe2e0981",
  1249 => x"069d3880",
  1250 => x"ff539fb5",
  1251 => x"2dbe8008",
  1252 => x"75708405",
  1253 => x"570cff13",
  1254 => x"53728025",
  1255 => x"ed388156",
  1256 => x"a7a904ff",
  1257 => x"145473c9",
  1258 => x"3881ff0b",
  1259 => x"d40c81ff",
  1260 => x"0bd40cd0",
  1261 => x"08708f2a",
  1262 => x"70810651",
  1263 => x"515372f3",
  1264 => x"3872d00c",
  1265 => x"75be800c",
  1266 => x"0298050d",
  1267 => x"0402f405",
  1268 => x"0d747088",
  1269 => x"2a83fe80",
  1270 => x"06707298",
  1271 => x"2a077288",
  1272 => x"2b87fc80",
  1273 => x"80067398",
  1274 => x"2b81f00a",
  1275 => x"06717307",
  1276 => x"07be800c",
  1277 => x"56515351",
  1278 => x"028c050d",
  1279 => x"0402f805",
  1280 => x"0d028e05",
  1281 => x"80f52d74",
  1282 => x"882b0770",
  1283 => x"83ffff06",
  1284 => x"be800c51",
  1285 => x"0288050d",
  1286 => x"0402fc05",
  1287 => x"0d725180",
  1288 => x"710c800b",
  1289 => x"84120c02",
  1290 => x"84050d04",
  1291 => x"02f0050d",
  1292 => x"75700884",
  1293 => x"12085353",
  1294 => x"53ff5471",
  1295 => x"712ea838",
  1296 => x"abf02d84",
  1297 => x"13087084",
  1298 => x"29148811",
  1299 => x"70087081",
  1300 => x"ff068418",
  1301 => x"08811187",
  1302 => x"06841a0c",
  1303 => x"53515551",
  1304 => x"5151abea",
  1305 => x"2d715473",
  1306 => x"be800c02",
  1307 => x"90050d04",
  1308 => x"02f8050d",
  1309 => x"abf02de0",
  1310 => x"08708b2a",
  1311 => x"70810651",
  1312 => x"52527080",
  1313 => x"2ea13880",
  1314 => x"c7f80870",
  1315 => x"842980c8",
  1316 => x"80057381",
  1317 => x"ff06710c",
  1318 => x"515180c7",
  1319 => x"f8088111",
  1320 => x"870680c7",
  1321 => x"f80c5180",
  1322 => x"0b80c8a0",
  1323 => x"0cabe32d",
  1324 => x"abea2d02",
  1325 => x"88050d04",
  1326 => x"02fc050d",
  1327 => x"abf02d81",
  1328 => x"0b80c8a0",
  1329 => x"0cabea2d",
  1330 => x"80c8a008",
  1331 => x"5170f938",
  1332 => x"0284050d",
  1333 => x"0402fc05",
  1334 => x"0d80c7f8",
  1335 => x"51a8992d",
  1336 => x"a8f051ab",
  1337 => x"df2dab89",
  1338 => x"2d028405",
  1339 => x"0d0402f4",
  1340 => x"050daaf0",
  1341 => x"04be8008",
  1342 => x"81f02e09",
  1343 => x"81068938",
  1344 => x"810bbdf4",
  1345 => x"0caaf004",
  1346 => x"be800881",
  1347 => x"e02e0981",
  1348 => x"06893881",
  1349 => x"0bbdf80c",
  1350 => x"aaf004be",
  1351 => x"800852bd",
  1352 => x"f808802e",
  1353 => x"8838be80",
  1354 => x"08818005",
  1355 => x"5271842c",
  1356 => x"728f0653",
  1357 => x"53bdf408",
  1358 => x"802e9938",
  1359 => x"728429bd",
  1360 => x"b4057213",
  1361 => x"81712b70",
  1362 => x"09730806",
  1363 => x"730c5153",
  1364 => x"53aae604",
  1365 => x"728429bd",
  1366 => x"b4057213",
  1367 => x"83712b72",
  1368 => x"0807720c",
  1369 => x"5353800b",
  1370 => x"bdf80c80",
  1371 => x"0bbdf40c",
  1372 => x"80c7f851",
  1373 => x"a8ac2dbe",
  1374 => x"8008ff24",
  1375 => x"fef73880",
  1376 => x"0bbe800c",
  1377 => x"028c050d",
  1378 => x"0402f805",
  1379 => x"0dbdb452",
  1380 => x"8f518072",
  1381 => x"70840554",
  1382 => x"0cff1151",
  1383 => x"708025f2",
  1384 => x"38028805",
  1385 => x"0d0402f0",
  1386 => x"050d7551",
  1387 => x"abf02d70",
  1388 => x"822cfc06",
  1389 => x"bdb41172",
  1390 => x"109e0671",
  1391 => x"0870722a",
  1392 => x"70830682",
  1393 => x"742b7009",
  1394 => x"7406760c",
  1395 => x"54515657",
  1396 => x"535153ab",
  1397 => x"ea2d71be",
  1398 => x"800c0290",
  1399 => x"050d0471",
  1400 => x"980c04ff",
  1401 => x"b008be80",
  1402 => x"0c04810b",
  1403 => x"ffb00c04",
  1404 => x"800bffb0",
  1405 => x"0c0402fc",
  1406 => x"050d810b",
  1407 => x"bdfc0c81",
  1408 => x"5184e62d",
  1409 => x"0284050d",
  1410 => x"0402fc05",
  1411 => x"0d800bbd",
  1412 => x"fc0c8051",
  1413 => x"84e62d02",
  1414 => x"84050d04",
  1415 => x"02ec050d",
  1416 => x"76548052",
  1417 => x"870b8815",
  1418 => x"80f52d56",
  1419 => x"53747224",
  1420 => x"8338a053",
  1421 => x"725182ef",
  1422 => x"2d81128b",
  1423 => x"1580f52d",
  1424 => x"54527272",
  1425 => x"25de3802",
  1426 => x"94050d04",
  1427 => x"02f0050d",
  1428 => x"80c8b008",
  1429 => x"5481f82d",
  1430 => x"800b80c8",
  1431 => x"b40c7308",
  1432 => x"802e8184",
  1433 => x"38820bbe",
  1434 => x"940c80c8",
  1435 => x"b4088f06",
  1436 => x"be900c73",
  1437 => x"08527183",
  1438 => x"2e963871",
  1439 => x"83268938",
  1440 => x"71812eaf",
  1441 => x"38add104",
  1442 => x"71852e9f",
  1443 => x"38add104",
  1444 => x"881480f5",
  1445 => x"2d841508",
  1446 => x"bac45354",
  1447 => x"5285f22d",
  1448 => x"71842913",
  1449 => x"70085252",
  1450 => x"add50473",
  1451 => x"51ac9c2d",
  1452 => x"add10480",
  1453 => x"c8a40888",
  1454 => x"15082c70",
  1455 => x"81065152",
  1456 => x"71802e87",
  1457 => x"38bac851",
  1458 => x"adce04ba",
  1459 => x"cc5185f2",
  1460 => x"2d841408",
  1461 => x"5185f22d",
  1462 => x"80c8b408",
  1463 => x"810580c8",
  1464 => x"b40c8c14",
  1465 => x"54acde04",
  1466 => x"0290050d",
  1467 => x"047180c8",
  1468 => x"b00caccc",
  1469 => x"2d80c8b4",
  1470 => x"08ff0580",
  1471 => x"c8b80c04",
  1472 => x"02e8050d",
  1473 => x"80c8b008",
  1474 => x"80c8bc08",
  1475 => x"575580f8",
  1476 => x"51aba62d",
  1477 => x"be800881",
  1478 => x"2a708106",
  1479 => x"5152719b",
  1480 => x"388751ab",
  1481 => x"a62dbe80",
  1482 => x"08812a70",
  1483 => x"81065152",
  1484 => x"71802eb1",
  1485 => x"38aebb04",
  1486 => x"a9ee2d87",
  1487 => x"51aba62d",
  1488 => x"be8008f4",
  1489 => x"38aecb04",
  1490 => x"a9ee2d80",
  1491 => x"f851aba6",
  1492 => x"2dbe8008",
  1493 => x"f338bdfc",
  1494 => x"08813270",
  1495 => x"bdfc0c70",
  1496 => x"525284e6",
  1497 => x"2d800b80",
  1498 => x"c8a80c80",
  1499 => x"0b80c8ac",
  1500 => x"0cbdfc08",
  1501 => x"82fd3880",
  1502 => x"da51aba6",
  1503 => x"2dbe8008",
  1504 => x"802e8c38",
  1505 => x"80c8a808",
  1506 => x"81800780",
  1507 => x"c8a80c80",
  1508 => x"d951aba6",
  1509 => x"2dbe8008",
  1510 => x"802e8c38",
  1511 => x"80c8a808",
  1512 => x"80c00780",
  1513 => x"c8a80c81",
  1514 => x"9451aba6",
  1515 => x"2dbe8008",
  1516 => x"802e8b38",
  1517 => x"80c8a808",
  1518 => x"900780c8",
  1519 => x"a80c8191",
  1520 => x"51aba62d",
  1521 => x"be800880",
  1522 => x"2e8b3880",
  1523 => x"c8a808a0",
  1524 => x"0780c8a8",
  1525 => x"0c81f551",
  1526 => x"aba62dbe",
  1527 => x"8008802e",
  1528 => x"8b3880c8",
  1529 => x"a8088107",
  1530 => x"80c8a80c",
  1531 => x"81f251ab",
  1532 => x"a62dbe80",
  1533 => x"08802e8b",
  1534 => x"3880c8a8",
  1535 => x"08820780",
  1536 => x"c8a80c81",
  1537 => x"eb51aba6",
  1538 => x"2dbe8008",
  1539 => x"802e8b38",
  1540 => x"80c8a808",
  1541 => x"840780c8",
  1542 => x"a80c81f4",
  1543 => x"51aba62d",
  1544 => x"be800880",
  1545 => x"2e8b3880",
  1546 => x"c8a80888",
  1547 => x"0780c8a8",
  1548 => x"0c80d851",
  1549 => x"aba62dbe",
  1550 => x"8008802e",
  1551 => x"8c3880c8",
  1552 => x"ac088180",
  1553 => x"0780c8ac",
  1554 => x"0c9251ab",
  1555 => x"a62dbe80",
  1556 => x"08802e8c",
  1557 => x"3880c8ac",
  1558 => x"0880c007",
  1559 => x"80c8ac0c",
  1560 => x"9451aba6",
  1561 => x"2dbe8008",
  1562 => x"802e8b38",
  1563 => x"80c8ac08",
  1564 => x"900780c8",
  1565 => x"ac0c9151",
  1566 => x"aba62dbe",
  1567 => x"8008802e",
  1568 => x"8b3880c8",
  1569 => x"ac08a007",
  1570 => x"80c8ac0c",
  1571 => x"9d51aba6",
  1572 => x"2dbe8008",
  1573 => x"802e8b38",
  1574 => x"80c8ac08",
  1575 => x"810780c8",
  1576 => x"ac0c9b51",
  1577 => x"aba62dbe",
  1578 => x"8008802e",
  1579 => x"8b3880c8",
  1580 => x"ac088207",
  1581 => x"80c8ac0c",
  1582 => x"9c51aba6",
  1583 => x"2dbe8008",
  1584 => x"802e8b38",
  1585 => x"80c8ac08",
  1586 => x"840780c8",
  1587 => x"ac0ca351",
  1588 => x"aba62dbe",
  1589 => x"8008802e",
  1590 => x"8b3880c8",
  1591 => x"ac088807",
  1592 => x"80c8ac0c",
  1593 => x"81fd51ab",
  1594 => x"a62d81fa",
  1595 => x"51aba62d",
  1596 => x"b7bb0481",
  1597 => x"f551aba6",
  1598 => x"2dbe8008",
  1599 => x"812a7081",
  1600 => x"06515271",
  1601 => x"802eb338",
  1602 => x"80c8b808",
  1603 => x"5271802e",
  1604 => x"8a38ff12",
  1605 => x"80c8b80c",
  1606 => x"b2ba0480",
  1607 => x"c8b40810",
  1608 => x"80c8b408",
  1609 => x"05708429",
  1610 => x"16515288",
  1611 => x"1208802e",
  1612 => x"8938ff51",
  1613 => x"88120852",
  1614 => x"712d81f2",
  1615 => x"51aba62d",
  1616 => x"be800881",
  1617 => x"2a708106",
  1618 => x"51527180",
  1619 => x"2eb43880",
  1620 => x"c8b408ff",
  1621 => x"1180c8b8",
  1622 => x"08565353",
  1623 => x"7372258a",
  1624 => x"38811480",
  1625 => x"c8b80cb3",
  1626 => x"82047210",
  1627 => x"13708429",
  1628 => x"16515288",
  1629 => x"1208802e",
  1630 => x"8938fe51",
  1631 => x"88120852",
  1632 => x"712d81fd",
  1633 => x"51aba62d",
  1634 => x"be800881",
  1635 => x"2a708106",
  1636 => x"51527180",
  1637 => x"2eb13880",
  1638 => x"c8b80880",
  1639 => x"2e8a3880",
  1640 => x"0b80c8b8",
  1641 => x"0cb3c704",
  1642 => x"80c8b408",
  1643 => x"1080c8b4",
  1644 => x"08057084",
  1645 => x"29165152",
  1646 => x"88120880",
  1647 => x"2e8938fd",
  1648 => x"51881208",
  1649 => x"52712d81",
  1650 => x"fa51aba6",
  1651 => x"2dbe8008",
  1652 => x"812a7081",
  1653 => x"06515271",
  1654 => x"802eb138",
  1655 => x"80c8b408",
  1656 => x"ff115452",
  1657 => x"80c8b808",
  1658 => x"73258938",
  1659 => x"7280c8b8",
  1660 => x"0cb48c04",
  1661 => x"71101270",
  1662 => x"84291651",
  1663 => x"52881208",
  1664 => x"802e8938",
  1665 => x"fc518812",
  1666 => x"0852712d",
  1667 => x"80c8b808",
  1668 => x"70535473",
  1669 => x"802e8a38",
  1670 => x"8c15ff15",
  1671 => x"5555b493",
  1672 => x"04820bbe",
  1673 => x"940c718f",
  1674 => x"06be900c",
  1675 => x"81eb51ab",
  1676 => x"a62dbe80",
  1677 => x"08812a70",
  1678 => x"81065152",
  1679 => x"71802ead",
  1680 => x"38740885",
  1681 => x"2e098106",
  1682 => x"a4388815",
  1683 => x"80f52dff",
  1684 => x"05527188",
  1685 => x"1681b72d",
  1686 => x"71982b52",
  1687 => x"71802588",
  1688 => x"38800b88",
  1689 => x"1681b72d",
  1690 => x"7451ac9c",
  1691 => x"2d81f451",
  1692 => x"aba62dbe",
  1693 => x"8008812a",
  1694 => x"70810651",
  1695 => x"5271802e",
  1696 => x"b3387408",
  1697 => x"852e0981",
  1698 => x"06aa3888",
  1699 => x"1580f52d",
  1700 => x"81055271",
  1701 => x"881681b7",
  1702 => x"2d7181ff",
  1703 => x"068b1680",
  1704 => x"f52d5452",
  1705 => x"72722787",
  1706 => x"38728816",
  1707 => x"81b72d74",
  1708 => x"51ac9c2d",
  1709 => x"80da51ab",
  1710 => x"a62dbe80",
  1711 => x"08812a70",
  1712 => x"81065152",
  1713 => x"71802e81",
  1714 => x"ac3880c8",
  1715 => x"b00880c8",
  1716 => x"b8085553",
  1717 => x"73802e8a",
  1718 => x"388c13ff",
  1719 => x"155553b5",
  1720 => x"d4047208",
  1721 => x"5271822e",
  1722 => x"a6387182",
  1723 => x"26893871",
  1724 => x"812eaa38",
  1725 => x"b6f50471",
  1726 => x"832eb438",
  1727 => x"71842e09",
  1728 => x"810680f1",
  1729 => x"38881308",
  1730 => x"51aded2d",
  1731 => x"b6f50480",
  1732 => x"c8b80851",
  1733 => x"88130852",
  1734 => x"712db6f5",
  1735 => x"04810b88",
  1736 => x"14082b80",
  1737 => x"c8a40832",
  1738 => x"80c8a40c",
  1739 => x"b6ca0488",
  1740 => x"1380f52d",
  1741 => x"81058b14",
  1742 => x"80f52d53",
  1743 => x"54717424",
  1744 => x"83388054",
  1745 => x"73881481",
  1746 => x"b72daccc",
  1747 => x"2db6f504",
  1748 => x"7508802e",
  1749 => x"a3387508",
  1750 => x"51aba62d",
  1751 => x"be800881",
  1752 => x"06527180",
  1753 => x"2e8c3880",
  1754 => x"c8b80851",
  1755 => x"84160852",
  1756 => x"712d8816",
  1757 => x"5675d938",
  1758 => x"8054800b",
  1759 => x"be940c73",
  1760 => x"8f06be90",
  1761 => x"0ca05273",
  1762 => x"80c8b808",
  1763 => x"2e098106",
  1764 => x"993880c8",
  1765 => x"b408ff05",
  1766 => x"74327009",
  1767 => x"81057072",
  1768 => x"079f2a91",
  1769 => x"71315151",
  1770 => x"53537151",
  1771 => x"82ef2d81",
  1772 => x"14548e74",
  1773 => x"25c438bd",
  1774 => x"fc085271",
  1775 => x"be800c02",
  1776 => x"98050d04",
  1777 => x"00ffffff",
  1778 => x"ff00ffff",
  1779 => x"ffff00ff",
  1780 => x"ffffff00",
  1781 => x"4f4b0000",
  1782 => x"52657365",
  1783 => x"74000000",
  1784 => x"53617665",
  1785 => x"20736574",
  1786 => x"74696e67",
  1787 => x"73000000",
  1788 => x"5363616e",
  1789 => x"6c696e65",
  1790 => x"73000000",
  1791 => x"4c6f6164",
  1792 => x"20524f4d",
  1793 => x"20100000",
  1794 => x"45786974",
  1795 => x"00000000",
  1796 => x"4a6f7973",
  1797 => x"7469636b",
  1798 => x"20737761",
  1799 => x"70000000",
  1800 => x"4a6f7973",
  1801 => x"7469636b",
  1802 => x"206e6f72",
  1803 => x"6d616c00",
  1804 => x"56474120",
  1805 => x"2d203331",
  1806 => x"4b487a2c",
  1807 => x"20363048",
  1808 => x"7a000000",
  1809 => x"5456202d",
  1810 => x"20343830",
  1811 => x"692c2036",
  1812 => x"30487a00",
  1813 => x"4261636b",
  1814 => x"00000000",
  1815 => x"4c6f6164",
  1816 => x"20457272",
  1817 => x"6f722100",
  1818 => x"46504741",
  1819 => x"47454e20",
  1820 => x"43464700",
  1821 => x"496e6974",
  1822 => x"69616c69",
  1823 => x"7a696e67",
  1824 => x"20534420",
  1825 => x"63617264",
  1826 => x"0a000000",
  1827 => x"424f4f54",
  1828 => x"20202020",
  1829 => x"47454e00",
  1830 => x"43617264",
  1831 => x"20696e69",
  1832 => x"74206661",
  1833 => x"696c6564",
  1834 => x"0a000000",
  1835 => x"4d425220",
  1836 => x"6661696c",
  1837 => x"0a000000",
  1838 => x"46415431",
  1839 => x"36202020",
  1840 => x"00000000",
  1841 => x"46415433",
  1842 => x"32202020",
  1843 => x"00000000",
  1844 => x"4e6f2070",
  1845 => x"61727469",
  1846 => x"74696f6e",
  1847 => x"20736967",
  1848 => x"0a000000",
  1849 => x"42616420",
  1850 => x"70617274",
  1851 => x"0a000000",
  1852 => x"53444843",
  1853 => x"20657272",
  1854 => x"6f72210a",
  1855 => x"00000000",
  1856 => x"53442069",
  1857 => x"6e69742e",
  1858 => x"2e2e0a00",
  1859 => x"53442063",
  1860 => x"61726420",
  1861 => x"72657365",
  1862 => x"74206661",
  1863 => x"696c6564",
  1864 => x"210a0000",
  1865 => x"57726974",
  1866 => x"65206661",
  1867 => x"696c6564",
  1868 => x"0a000000",
  1869 => x"52656164",
  1870 => x"20666169",
  1871 => x"6c65640a",
  1872 => x"00000000",
  1873 => x"16200000",
  1874 => x"14200000",
  1875 => x"15200000",
  1876 => x"00000002",
  1877 => x"00000000",
  1878 => x"00000002",
  1879 => x"00001bd8",
  1880 => x"000004aa",
  1881 => x"00000002",
  1882 => x"00001be0",
  1883 => x"0000037d",
  1884 => x"00000003",
  1885 => x"00001dc0",
  1886 => x"00000002",
  1887 => x"00000001",
  1888 => x"00001bf0",
  1889 => x"00000001",
  1890 => x"00000003",
  1891 => x"00001db8",
  1892 => x"00000002",
  1893 => x"00000002",
  1894 => x"00001bfc",
  1895 => x"00000759",
  1896 => x"00000002",
  1897 => x"00001c08",
  1898 => x"00001609",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00001c10",
  1903 => x"00001c20",
  1904 => x"00001c30",
  1905 => x"00001c44",
  1906 => x"00000002",
  1907 => x"00001f30",
  1908 => x"00000538",
  1909 => x"00000002",
  1910 => x"00001f4e",
  1911 => x"00000538",
  1912 => x"00000002",
  1913 => x"00001f6c",
  1914 => x"00000538",
  1915 => x"00000002",
  1916 => x"00001f8a",
  1917 => x"00000538",
  1918 => x"00000002",
  1919 => x"00001fa8",
  1920 => x"00000538",
  1921 => x"00000002",
  1922 => x"00001fc6",
  1923 => x"00000538",
  1924 => x"00000002",
  1925 => x"00001fe4",
  1926 => x"00000538",
  1927 => x"00000002",
  1928 => x"00002002",
  1929 => x"00000538",
  1930 => x"00000002",
  1931 => x"00002020",
  1932 => x"00000538",
  1933 => x"00000002",
  1934 => x"0000203e",
  1935 => x"00000538",
  1936 => x"00000002",
  1937 => x"0000205c",
  1938 => x"00000538",
  1939 => x"00000002",
  1940 => x"0000207a",
  1941 => x"00000538",
  1942 => x"00000002",
  1943 => x"00002098",
  1944 => x"00000538",
  1945 => x"00000004",
  1946 => x"00001c54",
  1947 => x"00001d58",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"000006ed",
  1951 => x"00000000",
  1952 => x"00000004",
  1953 => x"00001c5c",
  1954 => x"00001d58",
  1955 => x"00000004",
  1956 => x"00001cfc",
  1957 => x"00001d58",
  1958 => x"00000004",
  1959 => x"00001bd4",
  1960 => x"00001d58",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

