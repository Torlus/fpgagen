-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"f4080b0b",
    10 => x"0bbdf808",
    11 => x"0b0b0bbd",
    12 => x"fc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bdfc0c0b",
    16 => x"0b0bbdf8",
    17 => x"0c0b0b0b",
    18 => x"bdf40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb7e0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bdf47080",
    57 => x"c8b4278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518fce04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbe840c",
    65 => x"9f0bbe88",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"be8808ff",
    69 => x"05be880c",
    70 => x"be880880",
    71 => x"25eb38be",
    72 => x"8408ff05",
    73 => x"be840cbe",
    74 => x"84088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbe",
    94 => x"8408258f",
    95 => x"3882b32d",
    96 => x"be8408ff",
    97 => x"05be840c",
    98 => x"82f504be",
    99 => x"8408be88",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038be84",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"be880881",
   109 => x"05be880c",
   110 => x"be880851",
   111 => x"9f7125e2",
   112 => x"38800bbe",
   113 => x"880cbe84",
   114 => x"088105be",
   115 => x"840c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34be8808",
   120 => x"8105be88",
   121 => x"0cbe8808",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbe880c",
   125 => x"be840881",
   126 => x"05be840c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"be8c0cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbe",
   162 => x"8c0c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72be8c08",
   167 => x"8407be8c",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"bae00c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"be8c0852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c8980cba",
   200 => x"fc718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"bdf40c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b8f852be",
   211 => x"90519cb8",
   212 => x"2dbdf408",
   213 => x"802ea138",
   214 => x"80c1ac52",
   215 => x"be90519e",
   216 => x"f92d80c1",
   217 => x"ac08be9c",
   218 => x"0c80c1ac",
   219 => x"08fec00c",
   220 => x"80c1ac08",
   221 => x"5186932d",
   222 => x"0288050d",
   223 => x"0402f005",
   224 => x"0d805192",
   225 => x"872db8f8",
   226 => x"52be9051",
   227 => x"9cb82dbd",
   228 => x"f408802e",
   229 => x"a838be9c",
   230 => x"0880c1ac",
   231 => x"0c80c1b0",
   232 => x"5480fd53",
   233 => x"80747084",
   234 => x"05560cff",
   235 => x"13537280",
   236 => x"25f23880",
   237 => x"c1ac52be",
   238 => x"90519fa2",
   239 => x"2d029005",
   240 => x"0d0402d8",
   241 => x"050dbe9c",
   242 => x"08fec00c",
   243 => x"810bfec4",
   244 => x"0c840bfe",
   245 => x"c40c7b52",
   246 => x"be90519c",
   247 => x"b82dbdf4",
   248 => x"0853bdf4",
   249 => x"08802e81",
   250 => x"ba38be94",
   251 => x"0855800b",
   252 => x"ff165759",
   253 => x"75792e8b",
   254 => x"38811976",
   255 => x"812a5759",
   256 => x"75f738f7",
   257 => x"19759fff",
   258 => x"06545972",
   259 => x"802e8b38",
   260 => x"fc8015be",
   261 => x"9052559e",
   262 => x"cb2d74b0",
   263 => x"80802e09",
   264 => x"81068938",
   265 => x"820bfedc",
   266 => x"0c88c304",
   267 => x"74988080",
   268 => x"2e098106",
   269 => x"8938810b",
   270 => x"fedc0c88",
   271 => x"c304800b",
   272 => x"fedc0c81",
   273 => x"5a807525",
   274 => x"80d73878",
   275 => x"52755184",
   276 => x"812d80c1",
   277 => x"ac52be90",
   278 => x"519ef92d",
   279 => x"bdf40880",
   280 => x"2ea83880",
   281 => x"c1ac5883",
   282 => x"fc577770",
   283 => x"84055908",
   284 => x"7083ffff",
   285 => x"0671902a",
   286 => x"fec80cfe",
   287 => x"c80cfc18",
   288 => x"58537680",
   289 => x"25e43889",
   290 => x"9104bdf4",
   291 => x"085a8480",
   292 => x"55be9051",
   293 => x"9ecb2dfc",
   294 => x"80158117",
   295 => x"575588c5",
   296 => x"04795372",
   297 => x"bdf40c02",
   298 => x"a8050d04",
   299 => x"02fc050d",
   300 => x"ac9f2dfe",
   301 => x"c4518171",
   302 => x"0c82710c",
   303 => x"0284050d",
   304 => x"0402f405",
   305 => x"0d747678",
   306 => x"53545280",
   307 => x"71259738",
   308 => x"72708105",
   309 => x"5480f52d",
   310 => x"72708105",
   311 => x"5481b72d",
   312 => x"ff115170",
   313 => x"eb388072",
   314 => x"81b72d02",
   315 => x"8c050d04",
   316 => x"02e8050d",
   317 => x"77568070",
   318 => x"56547376",
   319 => x"24b33880",
   320 => x"c7bc0874",
   321 => x"2eab3873",
   322 => x"519a812d",
   323 => x"bdf408bd",
   324 => x"f4080981",
   325 => x"0570bdf4",
   326 => x"08079f2a",
   327 => x"77058117",
   328 => x"57575353",
   329 => x"74762489",
   330 => x"3880c7bc",
   331 => x"087426d7",
   332 => x"3872bdf4",
   333 => x"0c029805",
   334 => x"0d0402f4",
   335 => x"050dbda0",
   336 => x"08155189",
   337 => x"f02dbdf4",
   338 => x"08802e95",
   339 => x"388b53bd",
   340 => x"f4085280",
   341 => x"c5ac5189",
   342 => x"c12d80c5",
   343 => x"ac5187c2",
   344 => x"2dbae451",
   345 => x"ae832dac",
   346 => x"9f2d8051",
   347 => x"84e62d02",
   348 => x"8c050d04",
   349 => x"02dc050d",
   350 => x"80705a55",
   351 => x"74bda008",
   352 => x"25b13880",
   353 => x"c7bc0875",
   354 => x"2ea93878",
   355 => x"519a812d",
   356 => x"bdf40809",
   357 => x"810570bd",
   358 => x"f408079f",
   359 => x"2a760581",
   360 => x"1b5b5654",
   361 => x"74bda008",
   362 => x"25893880",
   363 => x"c7bc0879",
   364 => x"26d93880",
   365 => x"557880c7",
   366 => x"bc082781",
   367 => x"d0387851",
   368 => x"9a812dbd",
   369 => x"f408802e",
   370 => x"81a538bd",
   371 => x"f4088b05",
   372 => x"80f52d70",
   373 => x"842a7081",
   374 => x"06771078",
   375 => x"842b80c5",
   376 => x"ac0b80f5",
   377 => x"2d5c5c53",
   378 => x"51555673",
   379 => x"802e80c7",
   380 => x"38741682",
   381 => x"2b8db00b",
   382 => x"bbf4120c",
   383 => x"54777531",
   384 => x"10bea411",
   385 => x"55569074",
   386 => x"70810556",
   387 => x"81b72da0",
   388 => x"7481b72d",
   389 => x"7681ff06",
   390 => x"81165854",
   391 => x"73802e8a",
   392 => x"389c5380",
   393 => x"c5ac528c",
   394 => x"b0048b53",
   395 => x"bdf40852",
   396 => x"bea61651",
   397 => x"8ce70474",
   398 => x"16822b8a",
   399 => x"ba0bbbf4",
   400 => x"120c5476",
   401 => x"81ff0681",
   402 => x"16585473",
   403 => x"802e8a38",
   404 => x"9c5380c5",
   405 => x"ac528cdf",
   406 => x"048b53bd",
   407 => x"f4085277",
   408 => x"753110be",
   409 => x"a4055176",
   410 => x"5589c12d",
   411 => x"8d820474",
   412 => x"90297531",
   413 => x"7010bea4",
   414 => x"055154bd",
   415 => x"f4087481",
   416 => x"b72d8119",
   417 => x"59748b24",
   418 => x"a2388bb5",
   419 => x"04749029",
   420 => x"75317010",
   421 => x"bea4058c",
   422 => x"77315751",
   423 => x"54807481",
   424 => x"b72d9e14",
   425 => x"ff165654",
   426 => x"74f33802",
   427 => x"a4050d04",
   428 => x"02fc050d",
   429 => x"bda00813",
   430 => x"5189f02d",
   431 => x"bdf40880",
   432 => x"2e8838bd",
   433 => x"f4085192",
   434 => x"872d800b",
   435 => x"bda00c8a",
   436 => x"f42dace2",
   437 => x"2d028405",
   438 => x"0d0402fc",
   439 => x"050d7251",
   440 => x"70fd2ead",
   441 => x"3870fd24",
   442 => x"8a3870fc",
   443 => x"2e80c438",
   444 => x"8ebb0470",
   445 => x"fe2eb138",
   446 => x"70ff2e09",
   447 => x"8106bc38",
   448 => x"bda00851",
   449 => x"70802eb3",
   450 => x"38ff11bd",
   451 => x"a00c8ebb",
   452 => x"04bda008",
   453 => x"f00570bd",
   454 => x"a00c5170",
   455 => x"80259c38",
   456 => x"800bbda0",
   457 => x"0c8ebb04",
   458 => x"bda00881",
   459 => x"05bda00c",
   460 => x"8ebb04bd",
   461 => x"a0089005",
   462 => x"bda00c8a",
   463 => x"f42dace2",
   464 => x"2d028405",
   465 => x"0d0402fc",
   466 => x"050dbe9c",
   467 => x"08fb06be",
   468 => x"9c0c7251",
   469 => x"8aba2d02",
   470 => x"84050d04",
   471 => x"02fc050d",
   472 => x"be9c0884",
   473 => x"07be9c0c",
   474 => x"72518aba",
   475 => x"2d028405",
   476 => x"0d0402fc",
   477 => x"050d800b",
   478 => x"bda00c8a",
   479 => x"f42dbbec",
   480 => x"51ae832d",
   481 => x"bbd451ae",
   482 => x"962d0284",
   483 => x"050d0402",
   484 => x"f8050d80",
   485 => x"c8980882",
   486 => x"06bb840b",
   487 => x"80f52d52",
   488 => x"5270802e",
   489 => x"85387181",
   490 => x"0752bb9c",
   491 => x"0b80f52d",
   492 => x"5170802e",
   493 => x"85387184",
   494 => x"0752bea0",
   495 => x"08802e85",
   496 => x"38719007",
   497 => x"5271bdf4",
   498 => x"0c028805",
   499 => x"0d0402f4",
   500 => x"050d810b",
   501 => x"bea00c90",
   502 => x"5186932d",
   503 => x"a9eb2dac",
   504 => x"802da9ce",
   505 => x"2da9ce2d",
   506 => x"81f82d81",
   507 => x"5184e62d",
   508 => x"a9ce2da9",
   509 => x"ce2d8151",
   510 => x"84e62d81",
   511 => x"0bfec40c",
   512 => x"900bfec0",
   513 => x"0c840bfe",
   514 => x"c40c830b",
   515 => x"fecc0cb9",
   516 => x"845185f2",
   517 => x"2d8452a3",
   518 => x"d92d93a8",
   519 => x"2dbdf408",
   520 => x"802e8638",
   521 => x"fe5290b1",
   522 => x"04ff1252",
   523 => x"718024e7",
   524 => x"3871802e",
   525 => x"81833886",
   526 => x"c42db99c",
   527 => x"5187c22d",
   528 => x"bdf40880",
   529 => x"2e8f38ba",
   530 => x"e451ae83",
   531 => x"2d805184",
   532 => x"e62d90df",
   533 => x"04bdf408",
   534 => x"518ef22d",
   535 => x"ac8c2daa",
   536 => x"842dae9c",
   537 => x"2dbdf408",
   538 => x"80c89c08",
   539 => x"882b80c8",
   540 => x"a00807fe",
   541 => x"d80c538f",
   542 => x"8f2dbdf4",
   543 => x"08be9c08",
   544 => x"2ea238bd",
   545 => x"f408be9c",
   546 => x"0cbdf408",
   547 => x"fec00c84",
   548 => x"52725184",
   549 => x"e62da9ce",
   550 => x"2da9ce2d",
   551 => x"ff125271",
   552 => x"8025ee38",
   553 => x"72802e89",
   554 => x"388a0bfe",
   555 => x"c40c90df",
   556 => x"04820bfe",
   557 => x"c40c90df",
   558 => x"04b9a851",
   559 => x"85f22d80",
   560 => x"0bbdf40c",
   561 => x"028c050d",
   562 => x"0402e805",
   563 => x"0d77797b",
   564 => x"58555580",
   565 => x"53727625",
   566 => x"a3387470",
   567 => x"81055680",
   568 => x"f52d7470",
   569 => x"81055680",
   570 => x"f52d5252",
   571 => x"71712e86",
   572 => x"38815191",
   573 => x"fe048113",
   574 => x"5391d504",
   575 => x"805170bd",
   576 => x"f40c0298",
   577 => x"050d0402",
   578 => x"ec050d76",
   579 => x"5574802e",
   580 => x"be389a15",
   581 => x"80e02d51",
   582 => x"a8932dbd",
   583 => x"f408bdf4",
   584 => x"0880c7dc",
   585 => x"0cbdf408",
   586 => x"545480c7",
   587 => x"b808802e",
   588 => x"99389415",
   589 => x"80e02d51",
   590 => x"a8932dbd",
   591 => x"f408902b",
   592 => x"83fff00a",
   593 => x"06707507",
   594 => x"51537280",
   595 => x"c7dc0c80",
   596 => x"c7dc0853",
   597 => x"72802e9d",
   598 => x"3880c7b0",
   599 => x"08fe1471",
   600 => x"2980c7c4",
   601 => x"080580c7",
   602 => x"e00c7084",
   603 => x"2b80c7bc",
   604 => x"0c5493a3",
   605 => x"0480c7c8",
   606 => x"0880c7dc",
   607 => x"0c80c7cc",
   608 => x"0880c7e0",
   609 => x"0c80c7b8",
   610 => x"08802e8b",
   611 => x"3880c7b0",
   612 => x"08842b53",
   613 => x"939e0480",
   614 => x"c7d00884",
   615 => x"2b537280",
   616 => x"c7bc0c02",
   617 => x"94050d04",
   618 => x"02d8050d",
   619 => x"800b80c7",
   620 => x"b80c80c1",
   621 => x"ac528051",
   622 => x"a6c32dbd",
   623 => x"f40854bd",
   624 => x"f4088c38",
   625 => x"b9bc5185",
   626 => x"f22d7355",
   627 => x"99840480",
   628 => x"56810b80",
   629 => x"c7e40c88",
   630 => x"53b9c852",
   631 => x"80c1e251",
   632 => x"91c92dbd",
   633 => x"f408762e",
   634 => x"09810688",
   635 => x"38bdf408",
   636 => x"80c7e40c",
   637 => x"8853b9d4",
   638 => x"5280c1fe",
   639 => x"5191c92d",
   640 => x"bdf40888",
   641 => x"38bdf408",
   642 => x"80c7e40c",
   643 => x"80c7e408",
   644 => x"802e80fd",
   645 => x"3880c4f2",
   646 => x"0b80f52d",
   647 => x"80c4f30b",
   648 => x"80f52d71",
   649 => x"982b7190",
   650 => x"2b0780c4",
   651 => x"f40b80f5",
   652 => x"2d70882b",
   653 => x"720780c4",
   654 => x"f50b80f5",
   655 => x"2d710780",
   656 => x"c5aa0b80",
   657 => x"f52d80c5",
   658 => x"ab0b80f5",
   659 => x"2d71882b",
   660 => x"07535f54",
   661 => x"525a5657",
   662 => x"557381ab",
   663 => x"aa2e0981",
   664 => x"068d3875",
   665 => x"51a7e32d",
   666 => x"bdf40856",
   667 => x"94fc0473",
   668 => x"82d4d52e",
   669 => x"8738b9e0",
   670 => x"5195c104",
   671 => x"80c1ac52",
   672 => x"7551a6c3",
   673 => x"2dbdf408",
   674 => x"55bdf408",
   675 => x"802e83f4",
   676 => x"388853b9",
   677 => x"d45280c1",
   678 => x"fe5191c9",
   679 => x"2dbdf408",
   680 => x"8a38810b",
   681 => x"80c7b80c",
   682 => x"95c70488",
   683 => x"53b9c852",
   684 => x"80c1e251",
   685 => x"91c92dbd",
   686 => x"f408802e",
   687 => x"8a38b9f4",
   688 => x"5185f22d",
   689 => x"96a60480",
   690 => x"c5aa0b80",
   691 => x"f52d5473",
   692 => x"80d52e09",
   693 => x"810680ce",
   694 => x"3880c5ab",
   695 => x"0b80f52d",
   696 => x"547381aa",
   697 => x"2e098106",
   698 => x"bd38800b",
   699 => x"80c1ac0b",
   700 => x"80f52d56",
   701 => x"547481e9",
   702 => x"2e833881",
   703 => x"547481eb",
   704 => x"2e8c3880",
   705 => x"5573752e",
   706 => x"09810682",
   707 => x"f73880c1",
   708 => x"b70b80f5",
   709 => x"2d55748e",
   710 => x"3880c1b8",
   711 => x"0b80f52d",
   712 => x"5473822e",
   713 => x"86388055",
   714 => x"99840480",
   715 => x"c1b90b80",
   716 => x"f52d7080",
   717 => x"c7b00cff",
   718 => x"0580c7b4",
   719 => x"0c80c1ba",
   720 => x"0b80f52d",
   721 => x"80c1bb0b",
   722 => x"80f52d58",
   723 => x"76057782",
   724 => x"80290570",
   725 => x"80c7c00c",
   726 => x"80c1bc0b",
   727 => x"80f52d70",
   728 => x"80c7d40c",
   729 => x"80c7b808",
   730 => x"59575876",
   731 => x"802e81b5",
   732 => x"388853b9",
   733 => x"d45280c1",
   734 => x"fe5191c9",
   735 => x"2dbdf408",
   736 => x"82823880",
   737 => x"c7b00870",
   738 => x"842b80c7",
   739 => x"bc0c7080",
   740 => x"c7d00c80",
   741 => x"c1d10b80",
   742 => x"f52d80c1",
   743 => x"d00b80f5",
   744 => x"2d718280",
   745 => x"290580c1",
   746 => x"d20b80f5",
   747 => x"2d708480",
   748 => x"80291280",
   749 => x"c1d30b80",
   750 => x"f52d7081",
   751 => x"800a2912",
   752 => x"7080c7d8",
   753 => x"0c80c7d4",
   754 => x"08712980",
   755 => x"c7c00805",
   756 => x"7080c7c4",
   757 => x"0c80c1d9",
   758 => x"0b80f52d",
   759 => x"80c1d80b",
   760 => x"80f52d71",
   761 => x"82802905",
   762 => x"80c1da0b",
   763 => x"80f52d70",
   764 => x"84808029",
   765 => x"1280c1db",
   766 => x"0b80f52d",
   767 => x"70982b81",
   768 => x"f00a0672",
   769 => x"057080c7",
   770 => x"c80cfe11",
   771 => x"7e297705",
   772 => x"80c7cc0c",
   773 => x"52595243",
   774 => x"545e5152",
   775 => x"59525d57",
   776 => x"595798fd",
   777 => x"0480c1be",
   778 => x"0b80f52d",
   779 => x"80c1bd0b",
   780 => x"80f52d71",
   781 => x"82802905",
   782 => x"7080c7bc",
   783 => x"0c70a029",
   784 => x"83ff0570",
   785 => x"892a7080",
   786 => x"c7d00c80",
   787 => x"c1c30b80",
   788 => x"f52d80c1",
   789 => x"c20b80f5",
   790 => x"2d718280",
   791 => x"29057080",
   792 => x"c7d80c7b",
   793 => x"71291e70",
   794 => x"80c7cc0c",
   795 => x"7d80c7c8",
   796 => x"0c730580",
   797 => x"c7c40c55",
   798 => x"5e515155",
   799 => x"55805192",
   800 => x"872d8155",
   801 => x"74bdf40c",
   802 => x"02a8050d",
   803 => x"0402ec05",
   804 => x"0d767087",
   805 => x"2c7180ff",
   806 => x"06555654",
   807 => x"80c7b808",
   808 => x"8a387388",
   809 => x"2c7481ff",
   810 => x"06545580",
   811 => x"c1ac5280",
   812 => x"c7c00815",
   813 => x"51a6c32d",
   814 => x"bdf40854",
   815 => x"bdf40880",
   816 => x"2eb63880",
   817 => x"c7b80880",
   818 => x"2e993872",
   819 => x"842980c1",
   820 => x"ac057008",
   821 => x"5253a7e3",
   822 => x"2dbdf408",
   823 => x"f00a0653",
   824 => x"99f60472",
   825 => x"1080c1ac",
   826 => x"057080e0",
   827 => x"2d5253a8",
   828 => x"932dbdf4",
   829 => x"08537254",
   830 => x"73bdf40c",
   831 => x"0294050d",
   832 => x"0402e005",
   833 => x"0d797084",
   834 => x"2c80c7e0",
   835 => x"0805718f",
   836 => x"06525553",
   837 => x"728a3880",
   838 => x"c1ac5273",
   839 => x"51a6c32d",
   840 => x"72a02980",
   841 => x"c1ac0554",
   842 => x"807480f5",
   843 => x"2d565374",
   844 => x"732e8338",
   845 => x"81537481",
   846 => x"e52e81f1",
   847 => x"38817074",
   848 => x"06545872",
   849 => x"802e81e5",
   850 => x"388b1480",
   851 => x"f52d7083",
   852 => x"2a790658",
   853 => x"56769938",
   854 => x"bda40853",
   855 => x"72893872",
   856 => x"80c5ac0b",
   857 => x"81b72d76",
   858 => x"bda40c73",
   859 => x"539caf04",
   860 => x"758f2e09",
   861 => x"810681b5",
   862 => x"38749f06",
   863 => x"8d2980c5",
   864 => x"9f115153",
   865 => x"811480f5",
   866 => x"2d737081",
   867 => x"055581b7",
   868 => x"2d831480",
   869 => x"f52d7370",
   870 => x"81055581",
   871 => x"b72d8514",
   872 => x"80f52d73",
   873 => x"70810555",
   874 => x"81b72d87",
   875 => x"1480f52d",
   876 => x"73708105",
   877 => x"5581b72d",
   878 => x"891480f5",
   879 => x"2d737081",
   880 => x"055581b7",
   881 => x"2d8e1480",
   882 => x"f52d7370",
   883 => x"81055581",
   884 => x"b72d9014",
   885 => x"80f52d73",
   886 => x"70810555",
   887 => x"81b72d92",
   888 => x"1480f52d",
   889 => x"73708105",
   890 => x"5581b72d",
   891 => x"941480f5",
   892 => x"2d737081",
   893 => x"055581b7",
   894 => x"2d961480",
   895 => x"f52d7370",
   896 => x"81055581",
   897 => x"b72d9814",
   898 => x"80f52d73",
   899 => x"70810555",
   900 => x"81b72d9c",
   901 => x"1480f52d",
   902 => x"73708105",
   903 => x"5581b72d",
   904 => x"9e1480f5",
   905 => x"2d7381b7",
   906 => x"2d77bda4",
   907 => x"0c805372",
   908 => x"bdf40c02",
   909 => x"a0050d04",
   910 => x"02cc050d",
   911 => x"7e605e5a",
   912 => x"800b80c7",
   913 => x"dc0880c7",
   914 => x"e008595c",
   915 => x"56805880",
   916 => x"c7bc0878",
   917 => x"2e81b238",
   918 => x"778f06a0",
   919 => x"17575473",
   920 => x"913880c1",
   921 => x"ac527651",
   922 => x"811757a6",
   923 => x"c32d80c1",
   924 => x"ac568076",
   925 => x"80f52d56",
   926 => x"5474742e",
   927 => x"83388154",
   928 => x"7481e52e",
   929 => x"80f73881",
   930 => x"70750655",
   931 => x"5c73802e",
   932 => x"80eb388b",
   933 => x"1680f52d",
   934 => x"98065978",
   935 => x"80df388b",
   936 => x"537c5275",
   937 => x"5191c92d",
   938 => x"bdf40880",
   939 => x"d0389c16",
   940 => x"0851a7e3",
   941 => x"2dbdf408",
   942 => x"841b0c9a",
   943 => x"1680e02d",
   944 => x"51a8932d",
   945 => x"bdf408bd",
   946 => x"f408881c",
   947 => x"0cbdf408",
   948 => x"555580c7",
   949 => x"b808802e",
   950 => x"98389416",
   951 => x"80e02d51",
   952 => x"a8932dbd",
   953 => x"f408902b",
   954 => x"83fff00a",
   955 => x"06701651",
   956 => x"5473881b",
   957 => x"0c787a0c",
   958 => x"7b549ec2",
   959 => x"04811858",
   960 => x"80c7bc08",
   961 => x"7826fed0",
   962 => x"3880c7b8",
   963 => x"08802eb0",
   964 => x"387a5199",
   965 => x"8d2dbdf4",
   966 => x"08bdf408",
   967 => x"80ffffff",
   968 => x"f806555b",
   969 => x"7380ffff",
   970 => x"fff82e94",
   971 => x"38bdf408",
   972 => x"fe0580c7",
   973 => x"b0082980",
   974 => x"c7c40805",
   975 => x"579ccd04",
   976 => x"805473bd",
   977 => x"f40c02b4",
   978 => x"050d0402",
   979 => x"f4050d74",
   980 => x"70088105",
   981 => x"710c7008",
   982 => x"80c7b408",
   983 => x"06535371",
   984 => x"8e388813",
   985 => x"0851998d",
   986 => x"2dbdf408",
   987 => x"88140c81",
   988 => x"0bbdf40c",
   989 => x"028c050d",
   990 => x"0402f005",
   991 => x"0d758811",
   992 => x"08fe0580",
   993 => x"c7b00829",
   994 => x"80c7c408",
   995 => x"11720880",
   996 => x"c7b40806",
   997 => x"05795553",
   998 => x"5454a6c3",
   999 => x"2d029005",
  1000 => x"0d0402f0",
  1001 => x"050d7588",
  1002 => x"1108fe05",
  1003 => x"80c7b008",
  1004 => x"2980c7c4",
  1005 => x"08117208",
  1006 => x"80c7b408",
  1007 => x"06057955",
  1008 => x"535454a5",
  1009 => x"832d0290",
  1010 => x"050d0402",
  1011 => x"f4050dd4",
  1012 => x"5281ff72",
  1013 => x"0c710853",
  1014 => x"81ff720c",
  1015 => x"72882b83",
  1016 => x"fe800672",
  1017 => x"087081ff",
  1018 => x"06515253",
  1019 => x"81ff720c",
  1020 => x"72710788",
  1021 => x"2b720870",
  1022 => x"81ff0651",
  1023 => x"525381ff",
  1024 => x"720c7271",
  1025 => x"07882b72",
  1026 => x"087081ff",
  1027 => x"067207bd",
  1028 => x"f40c5253",
  1029 => x"028c050d",
  1030 => x"0402f405",
  1031 => x"0d747671",
  1032 => x"81ff06d4",
  1033 => x"0c535380",
  1034 => x"c7e80885",
  1035 => x"3871892b",
  1036 => x"5271982a",
  1037 => x"d40c7190",
  1038 => x"2a7081ff",
  1039 => x"06d40c51",
  1040 => x"71882a70",
  1041 => x"81ff06d4",
  1042 => x"0c517181",
  1043 => x"ff06d40c",
  1044 => x"72902a70",
  1045 => x"81ff06d4",
  1046 => x"0c51d408",
  1047 => x"7081ff06",
  1048 => x"515182b8",
  1049 => x"bf527081",
  1050 => x"ff2e0981",
  1051 => x"06943881",
  1052 => x"ff0bd40c",
  1053 => x"d4087081",
  1054 => x"ff06ff14",
  1055 => x"54515171",
  1056 => x"e53870bd",
  1057 => x"f40c028c",
  1058 => x"050d0402",
  1059 => x"fc050d81",
  1060 => x"c75181ff",
  1061 => x"0bd40cff",
  1062 => x"11517080",
  1063 => x"25f43802",
  1064 => x"84050d04",
  1065 => x"02f0050d",
  1066 => x"a18b2d8f",
  1067 => x"cf538052",
  1068 => x"87fc80f7",
  1069 => x"51a0992d",
  1070 => x"bdf40854",
  1071 => x"bdf40881",
  1072 => x"2e098106",
  1073 => x"a33881ff",
  1074 => x"0bd40c82",
  1075 => x"0a52849c",
  1076 => x"80e951a0",
  1077 => x"992dbdf4",
  1078 => x"088b3881",
  1079 => x"ff0bd40c",
  1080 => x"7353a1ee",
  1081 => x"04a18b2d",
  1082 => x"ff135372",
  1083 => x"c13872bd",
  1084 => x"f40c0290",
  1085 => x"050d0402",
  1086 => x"f4050d81",
  1087 => x"ff0bd40c",
  1088 => x"93538052",
  1089 => x"87fc80c1",
  1090 => x"51a0992d",
  1091 => x"bdf4088b",
  1092 => x"3881ff0b",
  1093 => x"d40c8153",
  1094 => x"a2a404a1",
  1095 => x"8b2dff13",
  1096 => x"5372df38",
  1097 => x"72bdf40c",
  1098 => x"028c050d",
  1099 => x"0402f005",
  1100 => x"0da18b2d",
  1101 => x"83aa5284",
  1102 => x"9c80c851",
  1103 => x"a0992dbd",
  1104 => x"f408812e",
  1105 => x"09810692",
  1106 => x"389fcb2d",
  1107 => x"bdf40883",
  1108 => x"ffff0653",
  1109 => x"7283aa2e",
  1110 => x"9738a1f7",
  1111 => x"2da2eb04",
  1112 => x"8154a3d0",
  1113 => x"04ba8051",
  1114 => x"85f22d80",
  1115 => x"54a3d004",
  1116 => x"81ff0bd4",
  1117 => x"0cb153a1",
  1118 => x"a42dbdf4",
  1119 => x"08802e80",
  1120 => x"c0388052",
  1121 => x"87fc80fa",
  1122 => x"51a0992d",
  1123 => x"bdf408b1",
  1124 => x"3881ff0b",
  1125 => x"d40cd408",
  1126 => x"5381ff0b",
  1127 => x"d40c81ff",
  1128 => x"0bd40c81",
  1129 => x"ff0bd40c",
  1130 => x"81ff0bd4",
  1131 => x"0c72862a",
  1132 => x"708106bd",
  1133 => x"f4085651",
  1134 => x"5372802e",
  1135 => x"9338a2e0",
  1136 => x"0472822e",
  1137 => x"ff9f38ff",
  1138 => x"135372ff",
  1139 => x"aa387254",
  1140 => x"73bdf40c",
  1141 => x"0290050d",
  1142 => x"0402f005",
  1143 => x"0d810b80",
  1144 => x"c7e80c84",
  1145 => x"54d00870",
  1146 => x"8f2a7081",
  1147 => x"06515153",
  1148 => x"72f33872",
  1149 => x"d00ca18b",
  1150 => x"2dba9051",
  1151 => x"85f22dd0",
  1152 => x"08708f2a",
  1153 => x"70810651",
  1154 => x"515372f3",
  1155 => x"38810bd0",
  1156 => x"0cb15380",
  1157 => x"5284d480",
  1158 => x"c051a099",
  1159 => x"2dbdf408",
  1160 => x"812ea138",
  1161 => x"72822e09",
  1162 => x"81068c38",
  1163 => x"ba9c5185",
  1164 => x"f22d8053",
  1165 => x"a4fa04ff",
  1166 => x"135372d7",
  1167 => x"38ff1454",
  1168 => x"73ffa238",
  1169 => x"a2ad2dbd",
  1170 => x"f40880c7",
  1171 => x"e80cbdf4",
  1172 => x"088b3881",
  1173 => x"5287fc80",
  1174 => x"d051a099",
  1175 => x"2d81ff0b",
  1176 => x"d40cd008",
  1177 => x"708f2a70",
  1178 => x"81065151",
  1179 => x"5372f338",
  1180 => x"72d00c81",
  1181 => x"ff0bd40c",
  1182 => x"815372bd",
  1183 => x"f40c0290",
  1184 => x"050d0402",
  1185 => x"e8050d78",
  1186 => x"5681ff0b",
  1187 => x"d40cd008",
  1188 => x"708f2a70",
  1189 => x"81065151",
  1190 => x"5372f338",
  1191 => x"82810bd0",
  1192 => x"0c81ff0b",
  1193 => x"d40c7752",
  1194 => x"87fc80d8",
  1195 => x"51a0992d",
  1196 => x"bdf40880",
  1197 => x"2e8c38ba",
  1198 => x"b45185f2",
  1199 => x"2d8153a6",
  1200 => x"ba0481ff",
  1201 => x"0bd40c81",
  1202 => x"fe0bd40c",
  1203 => x"80ff5575",
  1204 => x"70840557",
  1205 => x"0870982a",
  1206 => x"d40c7090",
  1207 => x"2c7081ff",
  1208 => x"06d40c54",
  1209 => x"70882c70",
  1210 => x"81ff06d4",
  1211 => x"0c547081",
  1212 => x"ff06d40c",
  1213 => x"54ff1555",
  1214 => x"748025d3",
  1215 => x"3881ff0b",
  1216 => x"d40c81ff",
  1217 => x"0bd40c81",
  1218 => x"ff0bd40c",
  1219 => x"868da054",
  1220 => x"81ff0bd4",
  1221 => x"0cd40881",
  1222 => x"ff065574",
  1223 => x"8738ff14",
  1224 => x"5473ed38",
  1225 => x"81ff0bd4",
  1226 => x"0cd00870",
  1227 => x"8f2a7081",
  1228 => x"06515153",
  1229 => x"72f33872",
  1230 => x"d00c72bd",
  1231 => x"f40c0298",
  1232 => x"050d0402",
  1233 => x"e8050d78",
  1234 => x"55805681",
  1235 => x"ff0bd40c",
  1236 => x"d008708f",
  1237 => x"2a708106",
  1238 => x"51515372",
  1239 => x"f3388281",
  1240 => x"0bd00c81",
  1241 => x"ff0bd40c",
  1242 => x"775287fc",
  1243 => x"80d151a0",
  1244 => x"992d80db",
  1245 => x"c6df54bd",
  1246 => x"f408802e",
  1247 => x"8a38bac4",
  1248 => x"5185f22d",
  1249 => x"a7da0481",
  1250 => x"ff0bd40c",
  1251 => x"d4087081",
  1252 => x"ff065153",
  1253 => x"7281fe2e",
  1254 => x"0981069d",
  1255 => x"3880ff53",
  1256 => x"9fcb2dbd",
  1257 => x"f4087570",
  1258 => x"8405570c",
  1259 => x"ff135372",
  1260 => x"8025ed38",
  1261 => x"8156a7bf",
  1262 => x"04ff1454",
  1263 => x"73c93881",
  1264 => x"ff0bd40c",
  1265 => x"81ff0bd4",
  1266 => x"0cd00870",
  1267 => x"8f2a7081",
  1268 => x"06515153",
  1269 => x"72f33872",
  1270 => x"d00c75bd",
  1271 => x"f40c0298",
  1272 => x"050d0402",
  1273 => x"f4050d74",
  1274 => x"70882a83",
  1275 => x"fe800670",
  1276 => x"72982a07",
  1277 => x"72882b87",
  1278 => x"fc808006",
  1279 => x"73982b81",
  1280 => x"f00a0671",
  1281 => x"730707bd",
  1282 => x"f40c5651",
  1283 => x"5351028c",
  1284 => x"050d0402",
  1285 => x"f8050d02",
  1286 => x"8e0580f5",
  1287 => x"2d74882b",
  1288 => x"077083ff",
  1289 => x"ff06bdf4",
  1290 => x"0c510288",
  1291 => x"050d0402",
  1292 => x"fc050d72",
  1293 => x"5180710c",
  1294 => x"800b8412",
  1295 => x"0c028405",
  1296 => x"0d0402f0",
  1297 => x"050d7570",
  1298 => x"08841208",
  1299 => x"535353ff",
  1300 => x"5471712e",
  1301 => x"a838ac86",
  1302 => x"2d841308",
  1303 => x"70842914",
  1304 => x"88117008",
  1305 => x"7081ff06",
  1306 => x"84180881",
  1307 => x"11870684",
  1308 => x"1a0c5351",
  1309 => x"55515151",
  1310 => x"ac802d71",
  1311 => x"5473bdf4",
  1312 => x"0c029005",
  1313 => x"0d0402f8",
  1314 => x"050dac86",
  1315 => x"2de00870",
  1316 => x"8b2a7081",
  1317 => x"06515252",
  1318 => x"70802ea1",
  1319 => x"3880c7ec",
  1320 => x"08708429",
  1321 => x"80c7f405",
  1322 => x"7381ff06",
  1323 => x"710c5151",
  1324 => x"80c7ec08",
  1325 => x"81118706",
  1326 => x"80c7ec0c",
  1327 => x"51800b80",
  1328 => x"c8940cab",
  1329 => x"f92dac80",
  1330 => x"2d028805",
  1331 => x"0d0402fc",
  1332 => x"050dac86",
  1333 => x"2d810b80",
  1334 => x"c8940cac",
  1335 => x"802d80c8",
  1336 => x"94085170",
  1337 => x"f9380284",
  1338 => x"050d0402",
  1339 => x"fc050d80",
  1340 => x"c7ec51a8",
  1341 => x"af2da986",
  1342 => x"51abf52d",
  1343 => x"ab9f2d02",
  1344 => x"84050d04",
  1345 => x"02f4050d",
  1346 => x"ab8604bd",
  1347 => x"f40881f0",
  1348 => x"2e098106",
  1349 => x"8938810b",
  1350 => x"bde80cab",
  1351 => x"8604bdf4",
  1352 => x"0881e02e",
  1353 => x"09810689",
  1354 => x"38810bbd",
  1355 => x"ec0cab86",
  1356 => x"04bdf408",
  1357 => x"52bdec08",
  1358 => x"802e8838",
  1359 => x"bdf40881",
  1360 => x"80055271",
  1361 => x"842c728f",
  1362 => x"065353bd",
  1363 => x"e808802e",
  1364 => x"99387284",
  1365 => x"29bda805",
  1366 => x"72138171",
  1367 => x"2b700973",
  1368 => x"0806730c",
  1369 => x"515353aa",
  1370 => x"fc047284",
  1371 => x"29bda805",
  1372 => x"72138371",
  1373 => x"2b720807",
  1374 => x"720c5353",
  1375 => x"800bbdec",
  1376 => x"0c800bbd",
  1377 => x"e80c80c7",
  1378 => x"ec51a8c2",
  1379 => x"2dbdf408",
  1380 => x"ff24fef7",
  1381 => x"38800bbd",
  1382 => x"f40c028c",
  1383 => x"050d0402",
  1384 => x"f8050dbd",
  1385 => x"a8528f51",
  1386 => x"80727084",
  1387 => x"05540cff",
  1388 => x"11517080",
  1389 => x"25f23802",
  1390 => x"88050d04",
  1391 => x"02f0050d",
  1392 => x"7551ac86",
  1393 => x"2d70822c",
  1394 => x"fc06bda8",
  1395 => x"1172109e",
  1396 => x"06710870",
  1397 => x"722a7083",
  1398 => x"0682742b",
  1399 => x"70097406",
  1400 => x"760c5451",
  1401 => x"56575351",
  1402 => x"53ac802d",
  1403 => x"71bdf40c",
  1404 => x"0290050d",
  1405 => x"0471980c",
  1406 => x"04ffb008",
  1407 => x"bdf40c04",
  1408 => x"810bffb0",
  1409 => x"0c04800b",
  1410 => x"ffb00c04",
  1411 => x"02fc050d",
  1412 => x"810bbdf0",
  1413 => x"0c815184",
  1414 => x"e62d0284",
  1415 => x"050d0402",
  1416 => x"fc050d80",
  1417 => x"0bbdf00c",
  1418 => x"805184e6",
  1419 => x"2d028405",
  1420 => x"0d0402ec",
  1421 => x"050d7654",
  1422 => x"8052870b",
  1423 => x"881580f5",
  1424 => x"2d565374",
  1425 => x"72248338",
  1426 => x"a0537251",
  1427 => x"82ef2d81",
  1428 => x"128b1580",
  1429 => x"f52d5452",
  1430 => x"727225de",
  1431 => x"38029405",
  1432 => x"0d0402f0",
  1433 => x"050d80c8",
  1434 => x"a4085481",
  1435 => x"f82d800b",
  1436 => x"80c8a80c",
  1437 => x"7308802e",
  1438 => x"81843882",
  1439 => x"0bbe880c",
  1440 => x"80c8a808",
  1441 => x"8f06be84",
  1442 => x"0c730852",
  1443 => x"71832e96",
  1444 => x"38718326",
  1445 => x"89387181",
  1446 => x"2eaf38ad",
  1447 => x"e7047185",
  1448 => x"2e9f38ad",
  1449 => x"e7048814",
  1450 => x"80f52d84",
  1451 => x"1508bad4",
  1452 => x"53545285",
  1453 => x"f22d7184",
  1454 => x"29137008",
  1455 => x"5252adeb",
  1456 => x"047351ac",
  1457 => x"b22dade7",
  1458 => x"0480c898",
  1459 => x"08881508",
  1460 => x"2c708106",
  1461 => x"51527180",
  1462 => x"2e8738ba",
  1463 => x"d851ade4",
  1464 => x"04badc51",
  1465 => x"85f22d84",
  1466 => x"14085185",
  1467 => x"f22d80c8",
  1468 => x"a8088105",
  1469 => x"80c8a80c",
  1470 => x"8c1454ac",
  1471 => x"f4040290",
  1472 => x"050d0471",
  1473 => x"80c8a40c",
  1474 => x"ace22d80",
  1475 => x"c8a808ff",
  1476 => x"0580c8ac",
  1477 => x"0c047180",
  1478 => x"c8b00c04",
  1479 => x"02e8050d",
  1480 => x"80c8a408",
  1481 => x"80c8b008",
  1482 => x"575580f8",
  1483 => x"51abbc2d",
  1484 => x"bdf40881",
  1485 => x"2a708106",
  1486 => x"5152719b",
  1487 => x"388751ab",
  1488 => x"bc2dbdf4",
  1489 => x"08812a70",
  1490 => x"81065152",
  1491 => x"71802eb1",
  1492 => x"38aed704",
  1493 => x"aa842d87",
  1494 => x"51abbc2d",
  1495 => x"bdf408f4",
  1496 => x"38aee704",
  1497 => x"aa842d80",
  1498 => x"f851abbc",
  1499 => x"2dbdf408",
  1500 => x"f338bdf0",
  1501 => x"08813270",
  1502 => x"bdf00c70",
  1503 => x"525284e6",
  1504 => x"2d800b80",
  1505 => x"c89c0c80",
  1506 => x"0b80c8a0",
  1507 => x"0cbdf008",
  1508 => x"82fd3880",
  1509 => x"da51abbc",
  1510 => x"2dbdf408",
  1511 => x"802e8c38",
  1512 => x"80c89c08",
  1513 => x"81800780",
  1514 => x"c89c0c80",
  1515 => x"d951abbc",
  1516 => x"2dbdf408",
  1517 => x"802e8c38",
  1518 => x"80c89c08",
  1519 => x"80c00780",
  1520 => x"c89c0c81",
  1521 => x"9451abbc",
  1522 => x"2dbdf408",
  1523 => x"802e8b38",
  1524 => x"80c89c08",
  1525 => x"900780c8",
  1526 => x"9c0c8191",
  1527 => x"51abbc2d",
  1528 => x"bdf40880",
  1529 => x"2e8b3880",
  1530 => x"c89c08a0",
  1531 => x"0780c89c",
  1532 => x"0c81f551",
  1533 => x"abbc2dbd",
  1534 => x"f408802e",
  1535 => x"8b3880c8",
  1536 => x"9c088107",
  1537 => x"80c89c0c",
  1538 => x"81f251ab",
  1539 => x"bc2dbdf4",
  1540 => x"08802e8b",
  1541 => x"3880c89c",
  1542 => x"08820780",
  1543 => x"c89c0c81",
  1544 => x"eb51abbc",
  1545 => x"2dbdf408",
  1546 => x"802e8b38",
  1547 => x"80c89c08",
  1548 => x"840780c8",
  1549 => x"9c0c81f4",
  1550 => x"51abbc2d",
  1551 => x"bdf40880",
  1552 => x"2e8b3880",
  1553 => x"c89c0888",
  1554 => x"0780c89c",
  1555 => x"0c80d851",
  1556 => x"abbc2dbd",
  1557 => x"f408802e",
  1558 => x"8c3880c8",
  1559 => x"a0088180",
  1560 => x"0780c8a0",
  1561 => x"0c9251ab",
  1562 => x"bc2dbdf4",
  1563 => x"08802e8c",
  1564 => x"3880c8a0",
  1565 => x"0880c007",
  1566 => x"80c8a00c",
  1567 => x"9451abbc",
  1568 => x"2dbdf408",
  1569 => x"802e8b38",
  1570 => x"80c8a008",
  1571 => x"900780c8",
  1572 => x"a00c9151",
  1573 => x"abbc2dbd",
  1574 => x"f408802e",
  1575 => x"8b3880c8",
  1576 => x"a008a007",
  1577 => x"80c8a00c",
  1578 => x"9d51abbc",
  1579 => x"2dbdf408",
  1580 => x"802e8b38",
  1581 => x"80c8a008",
  1582 => x"810780c8",
  1583 => x"a00c9b51",
  1584 => x"abbc2dbd",
  1585 => x"f408802e",
  1586 => x"8b3880c8",
  1587 => x"a0088207",
  1588 => x"80c8a00c",
  1589 => x"9c51abbc",
  1590 => x"2dbdf408",
  1591 => x"802e8b38",
  1592 => x"80c8a008",
  1593 => x"840780c8",
  1594 => x"a00ca351",
  1595 => x"abbc2dbd",
  1596 => x"f408802e",
  1597 => x"8b3880c8",
  1598 => x"a0088807",
  1599 => x"80c8a00c",
  1600 => x"81fd51ab",
  1601 => x"bc2d81fa",
  1602 => x"51abbc2d",
  1603 => x"b7d70481",
  1604 => x"f551abbc",
  1605 => x"2dbdf408",
  1606 => x"812a7081",
  1607 => x"06515271",
  1608 => x"802eb338",
  1609 => x"80c8ac08",
  1610 => x"5271802e",
  1611 => x"8a38ff12",
  1612 => x"80c8ac0c",
  1613 => x"b2d60480",
  1614 => x"c8a80810",
  1615 => x"80c8a808",
  1616 => x"05708429",
  1617 => x"16515288",
  1618 => x"1208802e",
  1619 => x"8938ff51",
  1620 => x"88120852",
  1621 => x"712d81f2",
  1622 => x"51abbc2d",
  1623 => x"bdf40881",
  1624 => x"2a708106",
  1625 => x"51527180",
  1626 => x"2eb43880",
  1627 => x"c8a808ff",
  1628 => x"1180c8ac",
  1629 => x"08565353",
  1630 => x"7372258a",
  1631 => x"38811480",
  1632 => x"c8ac0cb3",
  1633 => x"9e047210",
  1634 => x"13708429",
  1635 => x"16515288",
  1636 => x"1208802e",
  1637 => x"8938fe51",
  1638 => x"88120852",
  1639 => x"712d81fd",
  1640 => x"51abbc2d",
  1641 => x"bdf40881",
  1642 => x"2a708106",
  1643 => x"51527180",
  1644 => x"2eb13880",
  1645 => x"c8ac0880",
  1646 => x"2e8a3880",
  1647 => x"0b80c8ac",
  1648 => x"0cb3e304",
  1649 => x"80c8a808",
  1650 => x"1080c8a8",
  1651 => x"08057084",
  1652 => x"29165152",
  1653 => x"88120880",
  1654 => x"2e8938fd",
  1655 => x"51881208",
  1656 => x"52712d81",
  1657 => x"fa51abbc",
  1658 => x"2dbdf408",
  1659 => x"812a7081",
  1660 => x"06515271",
  1661 => x"802eb138",
  1662 => x"80c8a808",
  1663 => x"ff115452",
  1664 => x"80c8ac08",
  1665 => x"73258938",
  1666 => x"7280c8ac",
  1667 => x"0cb4a804",
  1668 => x"71101270",
  1669 => x"84291651",
  1670 => x"52881208",
  1671 => x"802e8938",
  1672 => x"fc518812",
  1673 => x"0852712d",
  1674 => x"80c8ac08",
  1675 => x"70535473",
  1676 => x"802e8a38",
  1677 => x"8c15ff15",
  1678 => x"5555b4af",
  1679 => x"04820bbe",
  1680 => x"880c718f",
  1681 => x"06be840c",
  1682 => x"81eb51ab",
  1683 => x"bc2dbdf4",
  1684 => x"08812a70",
  1685 => x"81065152",
  1686 => x"71802ead",
  1687 => x"38740885",
  1688 => x"2e098106",
  1689 => x"a4388815",
  1690 => x"80f52dff",
  1691 => x"05527188",
  1692 => x"1681b72d",
  1693 => x"71982b52",
  1694 => x"71802588",
  1695 => x"38800b88",
  1696 => x"1681b72d",
  1697 => x"7451acb2",
  1698 => x"2d81f451",
  1699 => x"abbc2dbd",
  1700 => x"f408812a",
  1701 => x"70810651",
  1702 => x"5271802e",
  1703 => x"b3387408",
  1704 => x"852e0981",
  1705 => x"06aa3888",
  1706 => x"1580f52d",
  1707 => x"81055271",
  1708 => x"881681b7",
  1709 => x"2d7181ff",
  1710 => x"068b1680",
  1711 => x"f52d5452",
  1712 => x"72722787",
  1713 => x"38728816",
  1714 => x"81b72d74",
  1715 => x"51acb22d",
  1716 => x"80da51ab",
  1717 => x"bc2dbdf4",
  1718 => x"08812a70",
  1719 => x"81065152",
  1720 => x"71802e81",
  1721 => x"ac3880c8",
  1722 => x"a40880c8",
  1723 => x"ac085553",
  1724 => x"73802e8a",
  1725 => x"388c13ff",
  1726 => x"155553b5",
  1727 => x"f0047208",
  1728 => x"5271822e",
  1729 => x"a6387182",
  1730 => x"26893871",
  1731 => x"812eaa38",
  1732 => x"b7910471",
  1733 => x"832eb438",
  1734 => x"71842e09",
  1735 => x"810680f1",
  1736 => x"38881308",
  1737 => x"51ae832d",
  1738 => x"b7910480",
  1739 => x"c8ac0851",
  1740 => x"88130852",
  1741 => x"712db791",
  1742 => x"04810b88",
  1743 => x"14082b80",
  1744 => x"c8980832",
  1745 => x"80c8980c",
  1746 => x"b6e60488",
  1747 => x"1380f52d",
  1748 => x"81058b14",
  1749 => x"80f52d53",
  1750 => x"54717424",
  1751 => x"83388054",
  1752 => x"73881481",
  1753 => x"b72dace2",
  1754 => x"2db79104",
  1755 => x"7508802e",
  1756 => x"a3387508",
  1757 => x"51abbc2d",
  1758 => x"bdf40881",
  1759 => x"06527180",
  1760 => x"2e8c3880",
  1761 => x"c8ac0851",
  1762 => x"84160852",
  1763 => x"712d8816",
  1764 => x"5675d938",
  1765 => x"8054800b",
  1766 => x"be880c73",
  1767 => x"8f06be84",
  1768 => x"0ca05273",
  1769 => x"80c8ac08",
  1770 => x"2e098106",
  1771 => x"993880c8",
  1772 => x"a808ff05",
  1773 => x"74327009",
  1774 => x"81057072",
  1775 => x"079f2a91",
  1776 => x"71315151",
  1777 => x"53537151",
  1778 => x"82ef2d81",
  1779 => x"14548e74",
  1780 => x"25c438bd",
  1781 => x"f0085271",
  1782 => x"bdf40c02",
  1783 => x"98050d04",
  1784 => x"00ffffff",
  1785 => x"ff00ffff",
  1786 => x"ffff00ff",
  1787 => x"ffffff00",
  1788 => x"52657365",
  1789 => x"74000000",
  1790 => x"53617665",
  1791 => x"20736574",
  1792 => x"74696e67",
  1793 => x"73000000",
  1794 => x"5363616e",
  1795 => x"6c696e65",
  1796 => x"73000000",
  1797 => x"4c6f6164",
  1798 => x"20524f4d",
  1799 => x"20100000",
  1800 => x"45786974",
  1801 => x"00000000",
  1802 => x"50432045",
  1803 => x"6e67696e",
  1804 => x"65206d6f",
  1805 => x"64650000",
  1806 => x"54757262",
  1807 => x"6f677261",
  1808 => x"66782031",
  1809 => x"36206d6f",
  1810 => x"64650000",
  1811 => x"56474120",
  1812 => x"2d203331",
  1813 => x"4b487a2c",
  1814 => x"20363048",
  1815 => x"7a000000",
  1816 => x"5456202d",
  1817 => x"20343830",
  1818 => x"692c2036",
  1819 => x"30487a00",
  1820 => x"4261636b",
  1821 => x"00000000",
  1822 => x"46504741",
  1823 => x"50434520",
  1824 => x"43464700",
  1825 => x"496e6974",
  1826 => x"69616c69",
  1827 => x"7a696e67",
  1828 => x"20534420",
  1829 => x"63617264",
  1830 => x"0a000000",
  1831 => x"424f4f54",
  1832 => x"20202020",
  1833 => x"50434500",
  1834 => x"43617264",
  1835 => x"20696e69",
  1836 => x"74206661",
  1837 => x"696c6564",
  1838 => x"0a000000",
  1839 => x"4d425220",
  1840 => x"6661696c",
  1841 => x"0a000000",
  1842 => x"46415431",
  1843 => x"36202020",
  1844 => x"00000000",
  1845 => x"46415433",
  1846 => x"32202020",
  1847 => x"00000000",
  1848 => x"4e6f2070",
  1849 => x"61727469",
  1850 => x"74696f6e",
  1851 => x"20736967",
  1852 => x"0a000000",
  1853 => x"42616420",
  1854 => x"70617274",
  1855 => x"0a000000",
  1856 => x"53444843",
  1857 => x"20657272",
  1858 => x"6f72210a",
  1859 => x"00000000",
  1860 => x"53442069",
  1861 => x"6e69742e",
  1862 => x"2e2e0a00",
  1863 => x"53442063",
  1864 => x"61726420",
  1865 => x"72657365",
  1866 => x"74206661",
  1867 => x"696c6564",
  1868 => x"210a0000",
  1869 => x"57726974",
  1870 => x"65206661",
  1871 => x"696c6564",
  1872 => x"0a000000",
  1873 => x"52656164",
  1874 => x"20666169",
  1875 => x"6c65640a",
  1876 => x"00000000",
  1877 => x"16200000",
  1878 => x"14200000",
  1879 => x"15200000",
  1880 => x"00000002",
  1881 => x"00000002",
  1882 => x"00001bf0",
  1883 => x"000004ac",
  1884 => x"00000002",
  1885 => x"00001bf8",
  1886 => x"0000037d",
  1887 => x"00000003",
  1888 => x"00001dcc",
  1889 => x"00000002",
  1890 => x"00000001",
  1891 => x"00001c08",
  1892 => x"00000001",
  1893 => x"00000003",
  1894 => x"00001dc4",
  1895 => x"00000002",
  1896 => x"00000002",
  1897 => x"00001c14",
  1898 => x"00000772",
  1899 => x"00000002",
  1900 => x"00001c20",
  1901 => x"0000161f",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00001c28",
  1906 => x"00001c38",
  1907 => x"00001c4c",
  1908 => x"00001c60",
  1909 => x"0000004d",
  1910 => x"00000746",
  1911 => x"0000002c",
  1912 => x"0000075c",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000002",
  1916 => x"00001f24",
  1917 => x"0000053a",
  1918 => x"00000002",
  1919 => x"00001f42",
  1920 => x"0000053a",
  1921 => x"00000002",
  1922 => x"00001f60",
  1923 => x"0000053a",
  1924 => x"00000002",
  1925 => x"00001f7e",
  1926 => x"0000053a",
  1927 => x"00000002",
  1928 => x"00001f9c",
  1929 => x"0000053a",
  1930 => x"00000002",
  1931 => x"00001fba",
  1932 => x"0000053a",
  1933 => x"00000002",
  1934 => x"00001fd8",
  1935 => x"0000053a",
  1936 => x"00000002",
  1937 => x"00001ff6",
  1938 => x"0000053a",
  1939 => x"00000002",
  1940 => x"00002014",
  1941 => x"0000053a",
  1942 => x"00000002",
  1943 => x"00002032",
  1944 => x"0000053a",
  1945 => x"00000002",
  1946 => x"00002050",
  1947 => x"0000053a",
  1948 => x"00000002",
  1949 => x"0000206e",
  1950 => x"0000053a",
  1951 => x"00000002",
  1952 => x"0000208c",
  1953 => x"0000053a",
  1954 => x"00000004",
  1955 => x"00001c70",
  1956 => x"00001d64",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"000006da",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

