-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM1;

architecture arch of CtrlROM_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b80c2",
     9 => x"90080b0b",
    10 => x"80c29408",
    11 => x"0b0b80c2",
    12 => x"98080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c2980c0b",
    16 => x"0b80c294",
    17 => x"0c0b0b80",
    18 => x"c2900c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbaec",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c29070",
    57 => x"80ccd027",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5190eb",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c2",
    65 => x"a00c9f0b",
    66 => x"80c2a40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c2a408ff",
    70 => x"0580c2a4",
    71 => x"0c80c2a4",
    72 => x"088025e8",
    73 => x"3880c2a0",
    74 => x"08ff0580",
    75 => x"c2a00c80",
    76 => x"c2a00880",
    77 => x"25d03802",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"80c2a008",
    97 => x"25913882",
    98 => x"bc2d80c2",
    99 => x"a008ff05",
   100 => x"80c2a00c",
   101 => x"82fe0480",
   102 => x"c2a00880",
   103 => x"c2a40853",
   104 => x"51728a2e",
   105 => x"098106be",
   106 => x"38715171",
   107 => x"9f24a438",
   108 => x"80c2a008",
   109 => x"a02911f8",
   110 => x"80115151",
   111 => x"a0713480",
   112 => x"c2a40881",
   113 => x"0580c2a4",
   114 => x"0c80c2a4",
   115 => x"08519f71",
   116 => x"25de3880",
   117 => x"0b80c2a4",
   118 => x"0c80c2a0",
   119 => x"08810580",
   120 => x"c2a00c83",
   121 => x"fc0470a0",
   122 => x"2912f880",
   123 => x"11515172",
   124 => x"713480c2",
   125 => x"a4088105",
   126 => x"80c2a40c",
   127 => x"80c2a408",
   128 => x"a02e0981",
   129 => x"06913880",
   130 => x"0b80c2a4",
   131 => x"0c80c2a0",
   132 => x"08810580",
   133 => x"c2a00c02",
   134 => x"8c050d04",
   135 => x"02e8050d",
   136 => x"77795656",
   137 => x"880bfc16",
   138 => x"77712c8f",
   139 => x"06545254",
   140 => x"80537272",
   141 => x"25953871",
   142 => x"53fbe014",
   143 => x"51877134",
   144 => x"8114ff14",
   145 => x"545472f1",
   146 => x"387153f9",
   147 => x"1576712c",
   148 => x"87065351",
   149 => x"71802e8b",
   150 => x"38fbe014",
   151 => x"51717134",
   152 => x"81145472",
   153 => x"8e249538",
   154 => x"8f733153",
   155 => x"fbe01451",
   156 => x"a0713481",
   157 => x"14ff1454",
   158 => x"5472f138",
   159 => x"0298050d",
   160 => x"0402ec05",
   161 => x"0d800b80",
   162 => x"c2a80cf6",
   163 => x"8c08f690",
   164 => x"0871882c",
   165 => x"565481ff",
   166 => x"06527372",
   167 => x"25893871",
   168 => x"54820b80",
   169 => x"c2a80c72",
   170 => x"882c7381",
   171 => x"ff065455",
   172 => x"7473258d",
   173 => x"387280c2",
   174 => x"a8088407",
   175 => x"80c2a80c",
   176 => x"5573842b",
   177 => x"87e87125",
   178 => x"83713170",
   179 => x"0b0b0bbe",
   180 => x"ac0c8171",
   181 => x"2bf6880c",
   182 => x"fea413ff",
   183 => x"122c7888",
   184 => x"29ff9405",
   185 => x"70812c80",
   186 => x"c2a80852",
   187 => x"58525551",
   188 => x"52547680",
   189 => x"2e853870",
   190 => x"81075170",
   191 => x"f6940c71",
   192 => x"098105f6",
   193 => x"800c7209",
   194 => x"8105f684",
   195 => x"0c029405",
   196 => x"0d0402f4",
   197 => x"050d7453",
   198 => x"72708105",
   199 => x"5480f52d",
   200 => x"5271802e",
   201 => x"89387151",
   202 => x"82f82d86",
   203 => x"9804028c",
   204 => x"050d0402",
   205 => x"f4050d74",
   206 => x"70820680",
   207 => x"ccb40cbe",
   208 => x"cc718106",
   209 => x"53535370",
   210 => x"881381b7",
   211 => x"2d981273",
   212 => x"822a7081",
   213 => x"06515252",
   214 => x"70881381",
   215 => x"b72d9812",
   216 => x"73832a70",
   217 => x"81065152",
   218 => x"52708813",
   219 => x"81b72d72",
   220 => x"842a7081",
   221 => x"06515372",
   222 => x"941381b7",
   223 => x"2d7080c2",
   224 => x"900c028c",
   225 => x"050d0402",
   226 => x"f8050dbc",
   227 => x"c45280c2",
   228 => x"ac519ee6",
   229 => x"2d80c290",
   230 => x"08802ea3",
   231 => x"3880c5c8",
   232 => x"5280c2ac",
   233 => x"51a1b32d",
   234 => x"80c5c808",
   235 => x"80c2b80c",
   236 => x"80c5c808",
   237 => x"fec00c80",
   238 => x"c5c80851",
   239 => x"86b32d02",
   240 => x"88050d04",
   241 => x"02f0050d",
   242 => x"8051949a",
   243 => x"2dbcc452",
   244 => x"80c2ac51",
   245 => x"9ee62d80",
   246 => x"c2900880",
   247 => x"2eaa3880",
   248 => x"c2b80880",
   249 => x"c5c80c80",
   250 => x"c5cc5480",
   251 => x"fd538074",
   252 => x"70840556",
   253 => x"0cff1353",
   254 => x"728025f2",
   255 => x"3880c5c8",
   256 => x"5280c2ac",
   257 => x"51a1dc2d",
   258 => x"0290050d",
   259 => x"0402d805",
   260 => x"0d800bbe",
   261 => x"b00c80c2",
   262 => x"b808fec0",
   263 => x"0c810bfe",
   264 => x"c40c840b",
   265 => x"fec40c7b",
   266 => x"5280c2ac",
   267 => x"519ee62d",
   268 => x"80c29008",
   269 => x"5380c290",
   270 => x"08802e81",
   271 => x"b83880c2",
   272 => x"b0085580",
   273 => x"0bff1657",
   274 => x"5975792e",
   275 => x"8b388119",
   276 => x"76812a57",
   277 => x"5975f738",
   278 => x"f7195974",
   279 => x"b080802e",
   280 => x"09810689",
   281 => x"38820bfe",
   282 => x"dc0c8984",
   283 => x"04749880",
   284 => x"802e0981",
   285 => x"06893881",
   286 => x"0bfedc0c",
   287 => x"89840480",
   288 => x"0bfedc0c",
   289 => x"815a8075",
   290 => x"2580e338",
   291 => x"78527551",
   292 => x"849c2d80",
   293 => x"c5c85280",
   294 => x"c2ac51a1",
   295 => x"b32d80c2",
   296 => x"9008802e",
   297 => x"a83880c5",
   298 => x"c85883fc",
   299 => x"57777084",
   300 => x"05590870",
   301 => x"83ffff06",
   302 => x"71902afe",
   303 => x"c80cfec8",
   304 => x"0cfc1858",
   305 => x"53768025",
   306 => x"e43889d5",
   307 => x"0480c290",
   308 => x"085a8480",
   309 => x"5580c2ac",
   310 => x"51a1832d",
   311 => x"fc801581",
   312 => x"17575574",
   313 => x"8024ffa4",
   314 => x"3879802e",
   315 => x"8638820b",
   316 => x"beb00c79",
   317 => x"537280c2",
   318 => x"900c02a8",
   319 => x"050d0402",
   320 => x"fc050daf",
   321 => x"872dfec4",
   322 => x"5181710c",
   323 => x"82710c02",
   324 => x"84050d04",
   325 => x"02f4050d",
   326 => x"74767853",
   327 => x"54528071",
   328 => x"25973872",
   329 => x"70810554",
   330 => x"80f52d72",
   331 => x"70810554",
   332 => x"81b72dff",
   333 => x"115170eb",
   334 => x"38807281",
   335 => x"b72d028c",
   336 => x"050d0402",
   337 => x"e8050d77",
   338 => x"56807056",
   339 => x"54737624",
   340 => x"b63880cb",
   341 => x"d808742e",
   342 => x"ae387351",
   343 => x"9cab2d80",
   344 => x"c2900880",
   345 => x"c2900809",
   346 => x"81057080",
   347 => x"c2900807",
   348 => x"9f2a7705",
   349 => x"81175757",
   350 => x"53537476",
   351 => x"24893880",
   352 => x"cbd80874",
   353 => x"26d43872",
   354 => x"80c2900c",
   355 => x"0298050d",
   356 => x"0402f405",
   357 => x"0d80c18c",
   358 => x"0815518a",
   359 => x"c32d80c2",
   360 => x"9008802e",
   361 => x"ac388b53",
   362 => x"80c29008",
   363 => x"5280c9c8",
   364 => x"518a942d",
   365 => x"80c9c851",
   366 => x"888d2d80",
   367 => x"c2900880",
   368 => x"2e8f38be",
   369 => x"b451b0ee",
   370 => x"2daf872d",
   371 => x"80518bdd",
   372 => x"0480c190",
   373 => x"51b0ee2d",
   374 => x"aef32d81",
   375 => x"5185812d",
   376 => x"028c050d",
   377 => x"0402dc05",
   378 => x"0d80705a",
   379 => x"557480c1",
   380 => x"8c0825b4",
   381 => x"3880cbd8",
   382 => x"08752eac",
   383 => x"3878519c",
   384 => x"ab2d80c2",
   385 => x"90080981",
   386 => x"057080c2",
   387 => x"9008079f",
   388 => x"2a760581",
   389 => x"1b5b5654",
   390 => x"7480c18c",
   391 => x"08258938",
   392 => x"80cbd808",
   393 => x"7926d638",
   394 => x"80557880",
   395 => x"cbd80827",
   396 => x"81d93878",
   397 => x"519cab2d",
   398 => x"80c29008",
   399 => x"802e81ab",
   400 => x"3880c290",
   401 => x"088b0580",
   402 => x"f52d7084",
   403 => x"2a708106",
   404 => x"77107884",
   405 => x"2b80c9c8",
   406 => x"0b80f52d",
   407 => x"5c5c5351",
   408 => x"55567380",
   409 => x"2e80ca38",
   410 => x"7416822b",
   411 => x"8eaf0bbf",
   412 => x"e0120c54",
   413 => x"77753110",
   414 => x"80c2c011",
   415 => x"55569074",
   416 => x"70810556",
   417 => x"81b72da0",
   418 => x"7481b72d",
   419 => x"7681ff06",
   420 => x"81165854",
   421 => x"73802e8a",
   422 => x"389c5380",
   423 => x"c9c8528d",
   424 => x"a9048b53",
   425 => x"80c29008",
   426 => x"5280c2c2",
   427 => x"16518de3",
   428 => x"04741682",
   429 => x"2b8b910b",
   430 => x"bfe0120c",
   431 => x"547681ff",
   432 => x"06811658",
   433 => x"5473802e",
   434 => x"8a389c53",
   435 => x"80c9c852",
   436 => x"8dda048b",
   437 => x"5380c290",
   438 => x"08527775",
   439 => x"311080c2",
   440 => x"c0055176",
   441 => x"558a942d",
   442 => x"8e800474",
   443 => x"90297531",
   444 => x"701080c2",
   445 => x"c0055154",
   446 => x"80c29008",
   447 => x"7481b72d",
   448 => x"81195974",
   449 => x"8b24a338",
   450 => x"8caa0474",
   451 => x"90297531",
   452 => x"701080c2",
   453 => x"c0058c77",
   454 => x"31575154",
   455 => x"807481b7",
   456 => x"2d9e14ff",
   457 => x"16565474",
   458 => x"f33802a4",
   459 => x"050d0402",
   460 => x"fc050d80",
   461 => x"c18c0813",
   462 => x"518ac32d",
   463 => x"80c29008",
   464 => x"802e8938",
   465 => x"80c29008",
   466 => x"51949a2d",
   467 => x"800b80c1",
   468 => x"8c0c8be5",
   469 => x"2dafcb2d",
   470 => x"0284050d",
   471 => x"0402fc05",
   472 => x"0d725170",
   473 => x"fd2eb038",
   474 => x"70fd248a",
   475 => x"3870fc2e",
   476 => x"80cc388f",
   477 => x"c80470fe",
   478 => x"2eb73870",
   479 => x"ff2e0981",
   480 => x"0680c538",
   481 => x"80c18c08",
   482 => x"5170802e",
   483 => x"bb38ff11",
   484 => x"80c18c0c",
   485 => x"8fc80480",
   486 => x"c18c08f0",
   487 => x"057080c1",
   488 => x"8c0c5170",
   489 => x"8025a138",
   490 => x"800b80c1",
   491 => x"8c0c8fc8",
   492 => x"0480c18c",
   493 => x"08810580",
   494 => x"c18c0c8f",
   495 => x"c80480c1",
   496 => x"8c089005",
   497 => x"80c18c0c",
   498 => x"8be52daf",
   499 => x"cb2d0284",
   500 => x"050d0402",
   501 => x"fc050d80",
   502 => x"0b80c18c",
   503 => x"0c8be52d",
   504 => x"bfd851b0",
   505 => x"ee2d0284",
   506 => x"050d04be",
   507 => x"f80b80f5",
   508 => x"2d80c290",
   509 => x"0c0402fc",
   510 => x"050d7287",
   511 => x"065170be",
   512 => x"f80b81b7",
   513 => x"2d028405",
   514 => x"0d0402f8",
   515 => x"050d80cc",
   516 => x"b4088206",
   517 => x"bed40b80",
   518 => x"f52d5252",
   519 => x"70802e85",
   520 => x"38718107",
   521 => x"52beec0b",
   522 => x"80f52d51",
   523 => x"70802e85",
   524 => x"38718407",
   525 => x"52bf840b",
   526 => x"80f52d51",
   527 => x"70802e85",
   528 => x"38718807",
   529 => x"52bf900b",
   530 => x"80f52d51",
   531 => x"70802e85",
   532 => x"38719007",
   533 => x"5280c2bc",
   534 => x"08802e85",
   535 => x"38719007",
   536 => x"527180c2",
   537 => x"900c0288",
   538 => x"050d0402",
   539 => x"f0050d81",
   540 => x"0b80c2bc",
   541 => x"0c800bbe",
   542 => x"b00c8753",
   543 => x"905186b3",
   544 => x"2d72518f",
   545 => x"f62d810b",
   546 => x"fec40c84",
   547 => x"0bfec40c",
   548 => x"830bfecc",
   549 => x"0cbcd051",
   550 => x"86922d84",
   551 => x"52a6a22d",
   552 => x"95c02d80",
   553 => x"c2900880",
   554 => x"2e8638fe",
   555 => x"5291b804",
   556 => x"ff125271",
   557 => x"8024e638",
   558 => x"71802e82",
   559 => x"8d38acc0",
   560 => x"2daee72d",
   561 => x"aca32dac",
   562 => x"a32d81f9",
   563 => x"2d815185",
   564 => x"812daca3",
   565 => x"2daca32d",
   566 => x"81518581",
   567 => x"2d87872d",
   568 => x"bce85188",
   569 => x"8d2d80c2",
   570 => x"9008802e",
   571 => x"9438beb4",
   572 => x"51b0ee2d",
   573 => x"80518581",
   574 => x"2d820bbe",
   575 => x"b00c928c",
   576 => x"0480c290",
   577 => x"08518fd3",
   578 => x"2daef32d",
   579 => x"acd92db1",
   580 => x"812d80c2",
   581 => x"900880cc",
   582 => x"b808882b",
   583 => x"80ccbc08",
   584 => x"07fed80c",
   585 => x"54908a2d",
   586 => x"80c29008",
   587 => x"80c2b808",
   588 => x"2ea53880",
   589 => x"c2900880",
   590 => x"c2b80c80",
   591 => x"c29008fe",
   592 => x"c00c8452",
   593 => x"73518581",
   594 => x"2daca32d",
   595 => x"aca32dff",
   596 => x"12527180",
   597 => x"25ee3885",
   598 => x"51aea02d",
   599 => x"80c29008",
   600 => x"812a7081",
   601 => x"06515271",
   602 => x"802e9538",
   603 => x"ff137009",
   604 => x"709f2c72",
   605 => x"06705452",
   606 => x"53538ff6",
   607 => x"2dafcb2d",
   608 => x"8651aea0",
   609 => x"2d80c290",
   610 => x"08812a70",
   611 => x"81065152",
   612 => x"71802e93",
   613 => x"38811353",
   614 => x"87732583",
   615 => x"38875372",
   616 => x"518ff62d",
   617 => x"afcb2d8f",
   618 => x"eb2d80c2",
   619 => x"9008fed4",
   620 => x"0c73802e",
   621 => x"8c38beb0",
   622 => x"088807fe",
   623 => x"c40c928c",
   624 => x"04beb008",
   625 => x"fec40c92",
   626 => x"8c04bcf4",
   627 => x"5186922d",
   628 => x"800b80c2",
   629 => x"900c0290",
   630 => x"050d0402",
   631 => x"e8050d77",
   632 => x"797b5855",
   633 => x"55805372",
   634 => x"7625a338",
   635 => x"74708105",
   636 => x"5680f52d",
   637 => x"74708105",
   638 => x"5680f52d",
   639 => x"52527171",
   640 => x"2e863881",
   641 => x"51949004",
   642 => x"81135393",
   643 => x"e7048051",
   644 => x"7080c290",
   645 => x"0c029805",
   646 => x"0d0402ec",
   647 => x"050d7655",
   648 => x"74802e80",
   649 => x"c2389a15",
   650 => x"80e02d51",
   651 => x"aae62d80",
   652 => x"c2900880",
   653 => x"c2900880",
   654 => x"cbf80c80",
   655 => x"c2900854",
   656 => x"5480cbd4",
   657 => x"08802e9a",
   658 => x"38941580",
   659 => x"e02d51aa",
   660 => x"e62d80c2",
   661 => x"9008902b",
   662 => x"83fff00a",
   663 => x"06707507",
   664 => x"51537280",
   665 => x"cbf80c80",
   666 => x"cbf80853",
   667 => x"72802e9d",
   668 => x"3880cbcc",
   669 => x"08fe1471",
   670 => x"2980cbe0",
   671 => x"080580cb",
   672 => x"fc0c7084",
   673 => x"2b80cbd8",
   674 => x"0c5495bb",
   675 => x"0480cbe4",
   676 => x"0880cbf8",
   677 => x"0c80cbe8",
   678 => x"0880cbfc",
   679 => x"0c80cbd4",
   680 => x"08802e8b",
   681 => x"3880cbcc",
   682 => x"08842b53",
   683 => x"95b60480",
   684 => x"cbec0884",
   685 => x"2b537280",
   686 => x"cbd80c02",
   687 => x"94050d04",
   688 => x"02d8050d",
   689 => x"800b80cb",
   690 => x"d40c80c5",
   691 => x"c8528051",
   692 => x"a9922d80",
   693 => x"c2900854",
   694 => x"80c29008",
   695 => x"8c38bd88",
   696 => x"5186922d",
   697 => x"73559ba8",
   698 => x"04805681",
   699 => x"0b80cc80",
   700 => x"0c8853bd",
   701 => x"945280c5",
   702 => x"fe5193db",
   703 => x"2d80c290",
   704 => x"08762e09",
   705 => x"81068938",
   706 => x"80c29008",
   707 => x"80cc800c",
   708 => x"8853bda0",
   709 => x"5280c69a",
   710 => x"5193db2d",
   711 => x"80c29008",
   712 => x"893880c2",
   713 => x"900880cc",
   714 => x"800c80cc",
   715 => x"8008802e",
   716 => x"81803880",
   717 => x"c98e0b80",
   718 => x"f52d80c9",
   719 => x"8f0b80f5",
   720 => x"2d71982b",
   721 => x"71902b07",
   722 => x"80c9900b",
   723 => x"80f52d70",
   724 => x"882b7207",
   725 => x"80c9910b",
   726 => x"80f52d71",
   727 => x"0780c9c6",
   728 => x"0b80f52d",
   729 => x"80c9c70b",
   730 => x"80f52d71",
   731 => x"882b0753",
   732 => x"5f54525a",
   733 => x"56575573",
   734 => x"81abaa2e",
   735 => x"0981068e",
   736 => x"387551aa",
   737 => x"b52d80c2",
   738 => x"90085697",
   739 => x"9b047382",
   740 => x"d4d52e87",
   741 => x"38bdac51",
   742 => x"97e40480",
   743 => x"c5c85275",
   744 => x"51a9922d",
   745 => x"80c29008",
   746 => x"5580c290",
   747 => x"08802e83",
   748 => x"f7388853",
   749 => x"bda05280",
   750 => x"c69a5193",
   751 => x"db2d80c2",
   752 => x"90088a38",
   753 => x"810b80cb",
   754 => x"d40c97ea",
   755 => x"048853bd",
   756 => x"945280c5",
   757 => x"fe5193db",
   758 => x"2d80c290",
   759 => x"08802e8a",
   760 => x"38bdc051",
   761 => x"86922d98",
   762 => x"c90480c9",
   763 => x"c60b80f5",
   764 => x"2d547380",
   765 => x"d52e0981",
   766 => x"0680ce38",
   767 => x"80c9c70b",
   768 => x"80f52d54",
   769 => x"7381aa2e",
   770 => x"098106bd",
   771 => x"38800b80",
   772 => x"c5c80b80",
   773 => x"f52d5654",
   774 => x"7481e92e",
   775 => x"83388154",
   776 => x"7481eb2e",
   777 => x"8c388055",
   778 => x"73752e09",
   779 => x"810682f8",
   780 => x"3880c5d3",
   781 => x"0b80f52d",
   782 => x"55748e38",
   783 => x"80c5d40b",
   784 => x"80f52d54",
   785 => x"73822e86",
   786 => x"3880559b",
   787 => x"a80480c5",
   788 => x"d50b80f5",
   789 => x"2d7080cb",
   790 => x"cc0cff05",
   791 => x"80cbd00c",
   792 => x"80c5d60b",
   793 => x"80f52d80",
   794 => x"c5d70b80",
   795 => x"f52d5876",
   796 => x"05778280",
   797 => x"29057080",
   798 => x"cbdc0c80",
   799 => x"c5d80b80",
   800 => x"f52d7080",
   801 => x"cbf00c80",
   802 => x"cbd40859",
   803 => x"57587680",
   804 => x"2e81b638",
   805 => x"8853bda0",
   806 => x"5280c69a",
   807 => x"5193db2d",
   808 => x"80c29008",
   809 => x"82823880",
   810 => x"cbcc0870",
   811 => x"842b80cb",
   812 => x"d80c7080",
   813 => x"cbec0c80",
   814 => x"c5ed0b80",
   815 => x"f52d80c5",
   816 => x"ec0b80f5",
   817 => x"2d718280",
   818 => x"290580c5",
   819 => x"ee0b80f5",
   820 => x"2d708480",
   821 => x"80291280",
   822 => x"c5ef0b80",
   823 => x"f52d7081",
   824 => x"800a2912",
   825 => x"7080cbf4",
   826 => x"0c80cbf0",
   827 => x"08712980",
   828 => x"cbdc0805",
   829 => x"7080cbe0",
   830 => x"0c80c5f5",
   831 => x"0b80f52d",
   832 => x"80c5f40b",
   833 => x"80f52d71",
   834 => x"82802905",
   835 => x"80c5f60b",
   836 => x"80f52d70",
   837 => x"84808029",
   838 => x"1280c5f7",
   839 => x"0b80f52d",
   840 => x"70982b81",
   841 => x"f00a0672",
   842 => x"057080cb",
   843 => x"e40cfe11",
   844 => x"7e297705",
   845 => x"80cbe80c",
   846 => x"52595243",
   847 => x"545e5152",
   848 => x"59525d57",
   849 => x"59579ba1",
   850 => x"0480c5da",
   851 => x"0b80f52d",
   852 => x"80c5d90b",
   853 => x"80f52d71",
   854 => x"82802905",
   855 => x"7080cbd8",
   856 => x"0c70a029",
   857 => x"83ff0570",
   858 => x"892a7080",
   859 => x"cbec0c80",
   860 => x"c5df0b80",
   861 => x"f52d80c5",
   862 => x"de0b80f5",
   863 => x"2d718280",
   864 => x"29057080",
   865 => x"cbf40c7b",
   866 => x"71291e70",
   867 => x"80cbe80c",
   868 => x"7d80cbe4",
   869 => x"0c730580",
   870 => x"cbe00c55",
   871 => x"5e515155",
   872 => x"55805194",
   873 => x"9a2d8155",
   874 => x"7480c290",
   875 => x"0c02a805",
   876 => x"0d0402ec",
   877 => x"050d7670",
   878 => x"872c7180",
   879 => x"ff065556",
   880 => x"5480cbd4",
   881 => x"088a3873",
   882 => x"882c7481",
   883 => x"ff065455",
   884 => x"80c5c852",
   885 => x"80cbdc08",
   886 => x"1551a992",
   887 => x"2d80c290",
   888 => x"085480c2",
   889 => x"9008802e",
   890 => x"b83880cb",
   891 => x"d408802e",
   892 => x"9a387284",
   893 => x"2980c5c8",
   894 => x"05700852",
   895 => x"53aab52d",
   896 => x"80c29008",
   897 => x"f00a0653",
   898 => x"9c9f0472",
   899 => x"1080c5c8",
   900 => x"057080e0",
   901 => x"2d5253aa",
   902 => x"e62d80c2",
   903 => x"90085372",
   904 => x"547380c2",
   905 => x"900c0294",
   906 => x"050d0402",
   907 => x"e0050d79",
   908 => x"70842c80",
   909 => x"cbfc0805",
   910 => x"718f0652",
   911 => x"5553728a",
   912 => x"3880c5c8",
   913 => x"527351a9",
   914 => x"922d72a0",
   915 => x"2980c5c8",
   916 => x"05548074",
   917 => x"80f52d56",
   918 => x"5374732e",
   919 => x"83388153",
   920 => x"7481e52e",
   921 => x"81f43881",
   922 => x"70740654",
   923 => x"5872802e",
   924 => x"81e8388b",
   925 => x"1480f52d",
   926 => x"70832a79",
   927 => x"06585676",
   928 => x"9b3880c1",
   929 => x"c0085372",
   930 => x"89387280",
   931 => x"c9c80b81",
   932 => x"b72d7680",
   933 => x"c1c00c73",
   934 => x"539edc04",
   935 => x"758f2e09",
   936 => x"810681b6",
   937 => x"38749f06",
   938 => x"8d2980c9",
   939 => x"bb115153",
   940 => x"811480f5",
   941 => x"2d737081",
   942 => x"055581b7",
   943 => x"2d831480",
   944 => x"f52d7370",
   945 => x"81055581",
   946 => x"b72d8514",
   947 => x"80f52d73",
   948 => x"70810555",
   949 => x"81b72d87",
   950 => x"1480f52d",
   951 => x"73708105",
   952 => x"5581b72d",
   953 => x"891480f5",
   954 => x"2d737081",
   955 => x"055581b7",
   956 => x"2d8e1480",
   957 => x"f52d7370",
   958 => x"81055581",
   959 => x"b72d9014",
   960 => x"80f52d73",
   961 => x"70810555",
   962 => x"81b72d92",
   963 => x"1480f52d",
   964 => x"73708105",
   965 => x"5581b72d",
   966 => x"941480f5",
   967 => x"2d737081",
   968 => x"055581b7",
   969 => x"2d961480",
   970 => x"f52d7370",
   971 => x"81055581",
   972 => x"b72d9814",
   973 => x"80f52d73",
   974 => x"70810555",
   975 => x"81b72d9c",
   976 => x"1480f52d",
   977 => x"73708105",
   978 => x"5581b72d",
   979 => x"9e1480f5",
   980 => x"2d7381b7",
   981 => x"2d7780c1",
   982 => x"c00c8053",
   983 => x"7280c290",
   984 => x"0c02a005",
   985 => x"0d0402cc",
   986 => x"050d7e60",
   987 => x"5e5a800b",
   988 => x"80cbf808",
   989 => x"80cbfc08",
   990 => x"595c5680",
   991 => x"5880cbd8",
   992 => x"08782e81",
   993 => x"b838778f",
   994 => x"06a01757",
   995 => x"54739138",
   996 => x"80c5c852",
   997 => x"76518117",
   998 => x"57a9922d",
   999 => x"80c5c856",
  1000 => x"807680f5",
  1001 => x"2d565474",
  1002 => x"742e8338",
  1003 => x"81547481",
  1004 => x"e52e80fd",
  1005 => x"38817075",
  1006 => x"06555c73",
  1007 => x"802e80f1",
  1008 => x"388b1680",
  1009 => x"f52d9806",
  1010 => x"597880e5",
  1011 => x"388b537c",
  1012 => x"52755193",
  1013 => x"db2d80c2",
  1014 => x"900880d5",
  1015 => x"389c1608",
  1016 => x"51aab52d",
  1017 => x"80c29008",
  1018 => x"841b0c9a",
  1019 => x"1680e02d",
  1020 => x"51aae62d",
  1021 => x"80c29008",
  1022 => x"80c29008",
  1023 => x"881c0c80",
  1024 => x"c2900855",
  1025 => x"5580cbd4",
  1026 => x"08802e99",
  1027 => x"38941680",
  1028 => x"e02d51aa",
  1029 => x"e62d80c2",
  1030 => x"9008902b",
  1031 => x"83fff00a",
  1032 => x"06701651",
  1033 => x"5473881b",
  1034 => x"0c787a0c",
  1035 => x"7b54a0f9",
  1036 => x"04811858",
  1037 => x"80cbd808",
  1038 => x"7826feca",
  1039 => x"3880cbd4",
  1040 => x"08802eb3",
  1041 => x"387a519b",
  1042 => x"b22d80c2",
  1043 => x"900880c2",
  1044 => x"900880ff",
  1045 => x"fffff806",
  1046 => x"555b7380",
  1047 => x"fffffff8",
  1048 => x"2e953880",
  1049 => x"c29008fe",
  1050 => x"0580cbcc",
  1051 => x"082980cb",
  1052 => x"e0080557",
  1053 => x"9efb0480",
  1054 => x"547380c2",
  1055 => x"900c02b4",
  1056 => x"050d0402",
  1057 => x"f4050d74",
  1058 => x"70088105",
  1059 => x"710c7008",
  1060 => x"80cbd008",
  1061 => x"06535371",
  1062 => x"8f388813",
  1063 => x"08519bb2",
  1064 => x"2d80c290",
  1065 => x"0888140c",
  1066 => x"810b80c2",
  1067 => x"900c028c",
  1068 => x"050d0402",
  1069 => x"f0050d75",
  1070 => x"881108fe",
  1071 => x"0580cbcc",
  1072 => x"082980cb",
  1073 => x"e0081172",
  1074 => x"0880cbd0",
  1075 => x"08060579",
  1076 => x"55535454",
  1077 => x"a9922d02",
  1078 => x"90050d04",
  1079 => x"02f0050d",
  1080 => x"75881108",
  1081 => x"fe0580cb",
  1082 => x"cc082980",
  1083 => x"cbe00811",
  1084 => x"720880cb",
  1085 => x"d0080605",
  1086 => x"79555354",
  1087 => x"54a7d02d",
  1088 => x"0290050d",
  1089 => x"0402f405",
  1090 => x"0dd45281",
  1091 => x"ff720c71",
  1092 => x"085381ff",
  1093 => x"720c7288",
  1094 => x"2b83fe80",
  1095 => x"06720870",
  1096 => x"81ff0651",
  1097 => x"525381ff",
  1098 => x"720c7271",
  1099 => x"07882b72",
  1100 => x"087081ff",
  1101 => x"06515253",
  1102 => x"81ff720c",
  1103 => x"72710788",
  1104 => x"2b720870",
  1105 => x"81ff0672",
  1106 => x"0780c290",
  1107 => x"0c525302",
  1108 => x"8c050d04",
  1109 => x"02f4050d",
  1110 => x"74767181",
  1111 => x"ff06d40c",
  1112 => x"535380cc",
  1113 => x"84088538",
  1114 => x"71892b52",
  1115 => x"71982ad4",
  1116 => x"0c71902a",
  1117 => x"7081ff06",
  1118 => x"d40c5171",
  1119 => x"882a7081",
  1120 => x"ff06d40c",
  1121 => x"517181ff",
  1122 => x"06d40c72",
  1123 => x"902a7081",
  1124 => x"ff06d40c",
  1125 => x"51d40870",
  1126 => x"81ff0651",
  1127 => x"5182b8bf",
  1128 => x"527081ff",
  1129 => x"2e098106",
  1130 => x"943881ff",
  1131 => x"0bd40cd4",
  1132 => x"087081ff",
  1133 => x"06ff1454",
  1134 => x"515171e5",
  1135 => x"387080c2",
  1136 => x"900c028c",
  1137 => x"050d0402",
  1138 => x"fc050d81",
  1139 => x"c75181ff",
  1140 => x"0bd40cff",
  1141 => x"11517080",
  1142 => x"25f43802",
  1143 => x"84050d04",
  1144 => x"02f0050d",
  1145 => x"a3c72d8f",
  1146 => x"cf538052",
  1147 => x"87fc80f7",
  1148 => x"51a2d42d",
  1149 => x"80c29008",
  1150 => x"5480c290",
  1151 => x"08812e09",
  1152 => x"8106a438",
  1153 => x"81ff0bd4",
  1154 => x"0c820a52",
  1155 => x"849c80e9",
  1156 => x"51a2d42d",
  1157 => x"80c29008",
  1158 => x"8b3881ff",
  1159 => x"0bd40c73",
  1160 => x"53a4ae04",
  1161 => x"a3c72dff",
  1162 => x"135372ff",
  1163 => x"bd387280",
  1164 => x"c2900c02",
  1165 => x"90050d04",
  1166 => x"02f4050d",
  1167 => x"81ff0bd4",
  1168 => x"0c935380",
  1169 => x"5287fc80",
  1170 => x"c151a2d4",
  1171 => x"2d80c290",
  1172 => x"088b3881",
  1173 => x"ff0bd40c",
  1174 => x"8153a4e6",
  1175 => x"04a3c72d",
  1176 => x"ff135372",
  1177 => x"de387280",
  1178 => x"c2900c02",
  1179 => x"8c050d04",
  1180 => x"02f0050d",
  1181 => x"a3c72d83",
  1182 => x"aa52849c",
  1183 => x"80c851a2",
  1184 => x"d42d80c2",
  1185 => x"9008812e",
  1186 => x"09810693",
  1187 => x"38a2852d",
  1188 => x"80c29008",
  1189 => x"83ffff06",
  1190 => x"537283aa",
  1191 => x"2e9738a4",
  1192 => x"b82da5b0",
  1193 => x"048154a6",
  1194 => x"9804bdcc",
  1195 => x"5186922d",
  1196 => x"8054a698",
  1197 => x"0481ff0b",
  1198 => x"d40cb153",
  1199 => x"a3e02d80",
  1200 => x"c2900880",
  1201 => x"2e80c238",
  1202 => x"805287fc",
  1203 => x"80fa51a2",
  1204 => x"d42d80c2",
  1205 => x"9008b238",
  1206 => x"81ff0bd4",
  1207 => x"0cd40853",
  1208 => x"81ff0bd4",
  1209 => x"0c81ff0b",
  1210 => x"d40c81ff",
  1211 => x"0bd40c81",
  1212 => x"ff0bd40c",
  1213 => x"72862a70",
  1214 => x"810680c2",
  1215 => x"90085651",
  1216 => x"5372802e",
  1217 => x"9338a5a5",
  1218 => x"0472822e",
  1219 => x"ff9c38ff",
  1220 => x"135372ff",
  1221 => x"a7387254",
  1222 => x"7380c290",
  1223 => x"0c029005",
  1224 => x"0d0402f0",
  1225 => x"050d810b",
  1226 => x"80cc840c",
  1227 => x"8454d008",
  1228 => x"708f2a70",
  1229 => x"81065151",
  1230 => x"5372f338",
  1231 => x"72d00ca3",
  1232 => x"c72dbddc",
  1233 => x"5186922d",
  1234 => x"d008708f",
  1235 => x"2a708106",
  1236 => x"51515372",
  1237 => x"f338810b",
  1238 => x"d00cb153",
  1239 => x"805284d4",
  1240 => x"80c051a2",
  1241 => x"d42d80c2",
  1242 => x"9008812e",
  1243 => x"a1387282",
  1244 => x"2e098106",
  1245 => x"8c38bde8",
  1246 => x"5186922d",
  1247 => x"8053a7c6",
  1248 => x"04ff1353",
  1249 => x"72d638ff",
  1250 => x"145473ff",
  1251 => x"a138a4f0",
  1252 => x"2d80c290",
  1253 => x"0880cc84",
  1254 => x"0c80c290",
  1255 => x"088b3881",
  1256 => x"5287fc80",
  1257 => x"d051a2d4",
  1258 => x"2d81ff0b",
  1259 => x"d40cd008",
  1260 => x"708f2a70",
  1261 => x"81065151",
  1262 => x"5372f338",
  1263 => x"72d00c81",
  1264 => x"ff0bd40c",
  1265 => x"81537280",
  1266 => x"c2900c02",
  1267 => x"90050d04",
  1268 => x"02e8050d",
  1269 => x"785681ff",
  1270 => x"0bd40cd0",
  1271 => x"08708f2a",
  1272 => x"70810651",
  1273 => x"515372f3",
  1274 => x"3882810b",
  1275 => x"d00c81ff",
  1276 => x"0bd40c77",
  1277 => x"5287fc80",
  1278 => x"d851a2d4",
  1279 => x"2d80c290",
  1280 => x"08802e8c",
  1281 => x"38be8051",
  1282 => x"86922d81",
  1283 => x"53a98804",
  1284 => x"81ff0bd4",
  1285 => x"0c81fe0b",
  1286 => x"d40c80ff",
  1287 => x"55757084",
  1288 => x"05570870",
  1289 => x"982ad40c",
  1290 => x"70902c70",
  1291 => x"81ff06d4",
  1292 => x"0c547088",
  1293 => x"2c7081ff",
  1294 => x"06d40c54",
  1295 => x"7081ff06",
  1296 => x"d40c54ff",
  1297 => x"15557480",
  1298 => x"25d33881",
  1299 => x"ff0bd40c",
  1300 => x"81ff0bd4",
  1301 => x"0c81ff0b",
  1302 => x"d40c868d",
  1303 => x"a05481ff",
  1304 => x"0bd40cd4",
  1305 => x"0881ff06",
  1306 => x"55748738",
  1307 => x"ff145473",
  1308 => x"ed3881ff",
  1309 => x"0bd40cd0",
  1310 => x"08708f2a",
  1311 => x"70810651",
  1312 => x"515372f3",
  1313 => x"3872d00c",
  1314 => x"7280c290",
  1315 => x"0c029805",
  1316 => x"0d0402e8",
  1317 => x"050d7855",
  1318 => x"805681ff",
  1319 => x"0bd40cd0",
  1320 => x"08708f2a",
  1321 => x"70810651",
  1322 => x"515372f3",
  1323 => x"3882810b",
  1324 => x"d00c81ff",
  1325 => x"0bd40c77",
  1326 => x"5287fc80",
  1327 => x"d151a2d4",
  1328 => x"2d80dbc6",
  1329 => x"df5480c2",
  1330 => x"9008802e",
  1331 => x"8a38be90",
  1332 => x"5186922d",
  1333 => x"aaab0481",
  1334 => x"ff0bd40c",
  1335 => x"d4087081",
  1336 => x"ff065153",
  1337 => x"7281fe2e",
  1338 => x"0981069e",
  1339 => x"3880ff53",
  1340 => x"a2852d80",
  1341 => x"c2900875",
  1342 => x"70840557",
  1343 => x"0cff1353",
  1344 => x"728025ec",
  1345 => x"388156aa",
  1346 => x"9004ff14",
  1347 => x"5473c838",
  1348 => x"81ff0bd4",
  1349 => x"0c81ff0b",
  1350 => x"d40cd008",
  1351 => x"708f2a70",
  1352 => x"81065151",
  1353 => x"5372f338",
  1354 => x"72d00c75",
  1355 => x"80c2900c",
  1356 => x"0298050d",
  1357 => x"0402f405",
  1358 => x"0d747088",
  1359 => x"2a83fe80",
  1360 => x"06707298",
  1361 => x"2a077288",
  1362 => x"2b87fc80",
  1363 => x"80067398",
  1364 => x"2b81f00a",
  1365 => x"06717307",
  1366 => x"0780c290",
  1367 => x"0c565153",
  1368 => x"51028c05",
  1369 => x"0d0402f8",
  1370 => x"050d028e",
  1371 => x"0580f52d",
  1372 => x"74882b07",
  1373 => x"7083ffff",
  1374 => x"0680c290",
  1375 => x"0c510288",
  1376 => x"050d0402",
  1377 => x"fc050d72",
  1378 => x"5180710c",
  1379 => x"800b8412",
  1380 => x"0c028405",
  1381 => x"0d0402f0",
  1382 => x"050d7570",
  1383 => x"08841208",
  1384 => x"535353ff",
  1385 => x"5471712e",
  1386 => x"a838aeed",
  1387 => x"2d841308",
  1388 => x"70842914",
  1389 => x"88117008",
  1390 => x"7081ff06",
  1391 => x"84180881",
  1392 => x"11870684",
  1393 => x"1a0c5351",
  1394 => x"55515151",
  1395 => x"aee72d71",
  1396 => x"547380c2",
  1397 => x"900c0290",
  1398 => x"050d0402",
  1399 => x"f8050dae",
  1400 => x"ed2de008",
  1401 => x"708b2a70",
  1402 => x"81065152",
  1403 => x"5270802e",
  1404 => x"a13880cc",
  1405 => x"88087084",
  1406 => x"2980cc90",
  1407 => x"057381ff",
  1408 => x"06710c51",
  1409 => x"5180cc88",
  1410 => x"08811187",
  1411 => x"0680cc88",
  1412 => x"0c51800b",
  1413 => x"80ccb00c",
  1414 => x"aedf2dae",
  1415 => x"e72d0288",
  1416 => x"050d0402",
  1417 => x"fc050dae",
  1418 => x"ed2d810b",
  1419 => x"80ccb00c",
  1420 => x"aee72d80",
  1421 => x"ccb00851",
  1422 => x"70f93802",
  1423 => x"84050d04",
  1424 => x"02fc050d",
  1425 => x"80cc8851",
  1426 => x"ab832dab",
  1427 => x"db51aedb",
  1428 => x"2dae822d",
  1429 => x"0284050d",
  1430 => x"0402f405",
  1431 => x"0dade704",
  1432 => x"80c29008",
  1433 => x"81f02e09",
  1434 => x"81068a38",
  1435 => x"810b80c2",
  1436 => x"840cade7",
  1437 => x"0480c290",
  1438 => x"0881e02e",
  1439 => x"0981068a",
  1440 => x"38810b80",
  1441 => x"c2880cad",
  1442 => x"e70480c2",
  1443 => x"90085280",
  1444 => x"c2880880",
  1445 => x"2e893880",
  1446 => x"c2900881",
  1447 => x"80055271",
  1448 => x"842c728f",
  1449 => x"06535380",
  1450 => x"c2840880",
  1451 => x"2e9a3872",
  1452 => x"842980c1",
  1453 => x"c4057213",
  1454 => x"81712b70",
  1455 => x"09730806",
  1456 => x"730c5153",
  1457 => x"53addb04",
  1458 => x"72842980",
  1459 => x"c1c40572",
  1460 => x"1383712b",
  1461 => x"72080772",
  1462 => x"0c535380",
  1463 => x"0b80c288",
  1464 => x"0c800b80",
  1465 => x"c2840c80",
  1466 => x"cc8851ab",
  1467 => x"962d80c2",
  1468 => x"9008ff24",
  1469 => x"feea3880",
  1470 => x"0b80c290",
  1471 => x"0c028c05",
  1472 => x"0d0402f8",
  1473 => x"050d80c1",
  1474 => x"c4528f51",
  1475 => x"80727084",
  1476 => x"05540cff",
  1477 => x"11517080",
  1478 => x"25f23802",
  1479 => x"88050d04",
  1480 => x"02f0050d",
  1481 => x"7551aeed",
  1482 => x"2d70822c",
  1483 => x"fc0680c1",
  1484 => x"c4117210",
  1485 => x"9e067108",
  1486 => x"70722a70",
  1487 => x"83068274",
  1488 => x"2b700974",
  1489 => x"06760c54",
  1490 => x"51565753",
  1491 => x"5153aee7",
  1492 => x"2d7180c2",
  1493 => x"900c0290",
  1494 => x"050d0471",
  1495 => x"980c04ff",
  1496 => x"b00880c2",
  1497 => x"900c0481",
  1498 => x"0bffb00c",
  1499 => x"04800bff",
  1500 => x"b00c0402",
  1501 => x"fc050d81",
  1502 => x"0b80c28c",
  1503 => x"0c815185",
  1504 => x"812d0284",
  1505 => x"050d0402",
  1506 => x"fc050d80",
  1507 => x"0b80c28c",
  1508 => x"0c805185",
  1509 => x"812d0284",
  1510 => x"050d0402",
  1511 => x"ec050d76",
  1512 => x"54805287",
  1513 => x"0b881580",
  1514 => x"f52d5653",
  1515 => x"74722483",
  1516 => x"38a05372",
  1517 => x"5182f82d",
  1518 => x"81128b15",
  1519 => x"80f52d54",
  1520 => x"52727225",
  1521 => x"de380294",
  1522 => x"050d0402",
  1523 => x"f0050d80",
  1524 => x"ccc00854",
  1525 => x"81f92d80",
  1526 => x"0b80ccc4",
  1527 => x"0c730880",
  1528 => x"2e818638",
  1529 => x"820b80c2",
  1530 => x"a40c80cc",
  1531 => x"c4088f06",
  1532 => x"80c2a00c",
  1533 => x"73085271",
  1534 => x"832e9638",
  1535 => x"71832689",
  1536 => x"3871812e",
  1537 => x"af38b0d2",
  1538 => x"0471852e",
  1539 => x"9f38b0d2",
  1540 => x"04881480",
  1541 => x"f52d8415",
  1542 => x"08bea053",
  1543 => x"54528692",
  1544 => x"2d718429",
  1545 => x"13700852",
  1546 => x"52b0d604",
  1547 => x"7351af9b",
  1548 => x"2db0d204",
  1549 => x"80ccb408",
  1550 => x"8815082c",
  1551 => x"70810651",
  1552 => x"5271802e",
  1553 => x"8738bea4",
  1554 => x"51b0cf04",
  1555 => x"bea85186",
  1556 => x"922d8414",
  1557 => x"08518692",
  1558 => x"2d80ccc4",
  1559 => x"08810580",
  1560 => x"ccc40c8c",
  1561 => x"1454afdd",
  1562 => x"04029005",
  1563 => x"0d047180",
  1564 => x"ccc00caf",
  1565 => x"cb2d80cc",
  1566 => x"c408ff05",
  1567 => x"80ccc80c",
  1568 => x"0402e805",
  1569 => x"0d80ccc0",
  1570 => x"0880cccc",
  1571 => x"08575580",
  1572 => x"f851aea0",
  1573 => x"2d80c290",
  1574 => x"08812a70",
  1575 => x"81065152",
  1576 => x"719c3887",
  1577 => x"51aea02d",
  1578 => x"80c29008",
  1579 => x"812a7081",
  1580 => x"06515271",
  1581 => x"802eb538",
  1582 => x"b1be04ac",
  1583 => x"d92d8751",
  1584 => x"aea02d80",
  1585 => x"c29008f3",
  1586 => x"38b1cf04",
  1587 => x"acd92d80",
  1588 => x"f851aea0",
  1589 => x"2d80c290",
  1590 => x"08f23880",
  1591 => x"c28c0881",
  1592 => x"327080c2",
  1593 => x"8c0c7052",
  1594 => x"5285812d",
  1595 => x"800b80cc",
  1596 => x"b80c800b",
  1597 => x"80ccbc0c",
  1598 => x"80c28c08",
  1599 => x"838d3880",
  1600 => x"da51aea0",
  1601 => x"2d80c290",
  1602 => x"08802e8c",
  1603 => x"3880ccb8",
  1604 => x"08818007",
  1605 => x"80ccb80c",
  1606 => x"80d951ae",
  1607 => x"a02d80c2",
  1608 => x"9008802e",
  1609 => x"8c3880cc",
  1610 => x"b80880c0",
  1611 => x"0780ccb8",
  1612 => x"0c819451",
  1613 => x"aea02d80",
  1614 => x"c2900880",
  1615 => x"2e8b3880",
  1616 => x"ccb80890",
  1617 => x"0780ccb8",
  1618 => x"0c819151",
  1619 => x"aea02d80",
  1620 => x"c2900880",
  1621 => x"2e8b3880",
  1622 => x"ccb808a0",
  1623 => x"0780ccb8",
  1624 => x"0c81f551",
  1625 => x"aea02d80",
  1626 => x"c2900880",
  1627 => x"2e8b3880",
  1628 => x"ccb80881",
  1629 => x"0780ccb8",
  1630 => x"0c81f251",
  1631 => x"aea02d80",
  1632 => x"c2900880",
  1633 => x"2e8b3880",
  1634 => x"ccb80882",
  1635 => x"0780ccb8",
  1636 => x"0c81eb51",
  1637 => x"aea02d80",
  1638 => x"c2900880",
  1639 => x"2e8b3880",
  1640 => x"ccb80884",
  1641 => x"0780ccb8",
  1642 => x"0c81f451",
  1643 => x"aea02d80",
  1644 => x"c2900880",
  1645 => x"2e8b3880",
  1646 => x"ccb80888",
  1647 => x"0780ccb8",
  1648 => x"0c80d851",
  1649 => x"aea02d80",
  1650 => x"c2900880",
  1651 => x"2e8c3880",
  1652 => x"ccbc0881",
  1653 => x"800780cc",
  1654 => x"bc0c9251",
  1655 => x"aea02d80",
  1656 => x"c2900880",
  1657 => x"2e8c3880",
  1658 => x"ccbc0880",
  1659 => x"c00780cc",
  1660 => x"bc0c9451",
  1661 => x"aea02d80",
  1662 => x"c2900880",
  1663 => x"2e8b3880",
  1664 => x"ccbc0890",
  1665 => x"0780ccbc",
  1666 => x"0c9151ae",
  1667 => x"a02d80c2",
  1668 => x"9008802e",
  1669 => x"8b3880cc",
  1670 => x"bc08a007",
  1671 => x"80ccbc0c",
  1672 => x"9d51aea0",
  1673 => x"2d80c290",
  1674 => x"08802e8b",
  1675 => x"3880ccbc",
  1676 => x"08810780",
  1677 => x"ccbc0c9b",
  1678 => x"51aea02d",
  1679 => x"80c29008",
  1680 => x"802e8b38",
  1681 => x"80ccbc08",
  1682 => x"820780cc",
  1683 => x"bc0c9c51",
  1684 => x"aea02d80",
  1685 => x"c2900880",
  1686 => x"2e8b3880",
  1687 => x"ccbc0884",
  1688 => x"0780ccbc",
  1689 => x"0ca351ae",
  1690 => x"a02d80c2",
  1691 => x"9008802e",
  1692 => x"8b3880cc",
  1693 => x"bc088807",
  1694 => x"80ccbc0c",
  1695 => x"81fd51ae",
  1696 => x"a02d81fa",
  1697 => x"51aea02d",
  1698 => x"bae00481",
  1699 => x"f551aea0",
  1700 => x"2d80c290",
  1701 => x"08812a70",
  1702 => x"81065152",
  1703 => x"71802eb3",
  1704 => x"3880ccc8",
  1705 => x"08527180",
  1706 => x"2e8a38ff",
  1707 => x"1280ccc8",
  1708 => x"0cb5d304",
  1709 => x"80ccc408",
  1710 => x"1080ccc4",
  1711 => x"08057084",
  1712 => x"29165152",
  1713 => x"88120880",
  1714 => x"2e8938ff",
  1715 => x"51881208",
  1716 => x"52712d81",
  1717 => x"f251aea0",
  1718 => x"2d80c290",
  1719 => x"08812a70",
  1720 => x"81065152",
  1721 => x"71802eb4",
  1722 => x"3880ccc4",
  1723 => x"08ff1180",
  1724 => x"ccc80856",
  1725 => x"53537372",
  1726 => x"258a3881",
  1727 => x"1480ccc8",
  1728 => x"0cb69c04",
  1729 => x"72101370",
  1730 => x"84291651",
  1731 => x"52881208",
  1732 => x"802e8938",
  1733 => x"fe518812",
  1734 => x"0852712d",
  1735 => x"81fd51ae",
  1736 => x"a02d80c2",
  1737 => x"9008812a",
  1738 => x"70810651",
  1739 => x"5271802e",
  1740 => x"b13880cc",
  1741 => x"c808802e",
  1742 => x"8a38800b",
  1743 => x"80ccc80c",
  1744 => x"b6e20480",
  1745 => x"ccc40810",
  1746 => x"80ccc408",
  1747 => x"05708429",
  1748 => x"16515288",
  1749 => x"1208802e",
  1750 => x"8938fd51",
  1751 => x"88120852",
  1752 => x"712d81fa",
  1753 => x"51aea02d",
  1754 => x"80c29008",
  1755 => x"812a7081",
  1756 => x"06515271",
  1757 => x"802eb138",
  1758 => x"80ccc408",
  1759 => x"ff115452",
  1760 => x"80ccc808",
  1761 => x"73258938",
  1762 => x"7280ccc8",
  1763 => x"0cb7a804",
  1764 => x"71101270",
  1765 => x"84291651",
  1766 => x"52881208",
  1767 => x"802e8938",
  1768 => x"fc518812",
  1769 => x"0852712d",
  1770 => x"80ccc808",
  1771 => x"70535473",
  1772 => x"802e8a38",
  1773 => x"8c15ff15",
  1774 => x"5555b7af",
  1775 => x"04820b80",
  1776 => x"c2a40c71",
  1777 => x"8f0680c2",
  1778 => x"a00c81eb",
  1779 => x"51aea02d",
  1780 => x"80c29008",
  1781 => x"812a7081",
  1782 => x"06515271",
  1783 => x"802ead38",
  1784 => x"7408852e",
  1785 => x"098106a4",
  1786 => x"38881580",
  1787 => x"f52dff05",
  1788 => x"52718816",
  1789 => x"81b72d71",
  1790 => x"982b5271",
  1791 => x"80258838",
  1792 => x"800b8816",
  1793 => x"81b72d74",
  1794 => x"51af9b2d",
  1795 => x"81f451ae",
  1796 => x"a02d80c2",
  1797 => x"9008812a",
  1798 => x"70810651",
  1799 => x"5271802e",
  1800 => x"b3387408",
  1801 => x"852e0981",
  1802 => x"06aa3888",
  1803 => x"1580f52d",
  1804 => x"81055271",
  1805 => x"881681b7",
  1806 => x"2d7181ff",
  1807 => x"068b1680",
  1808 => x"f52d5452",
  1809 => x"72722787",
  1810 => x"38728816",
  1811 => x"81b72d74",
  1812 => x"51af9b2d",
  1813 => x"80da51ae",
  1814 => x"a02d80c2",
  1815 => x"9008812a",
  1816 => x"70810651",
  1817 => x"5271802e",
  1818 => x"81ad3880",
  1819 => x"ccc00880",
  1820 => x"ccc80855",
  1821 => x"5373802e",
  1822 => x"8a388c13",
  1823 => x"ff155553",
  1824 => x"b8f50472",
  1825 => x"08527182",
  1826 => x"2ea63871",
  1827 => x"82268938",
  1828 => x"71812eaa",
  1829 => x"38ba9704",
  1830 => x"71832eb4",
  1831 => x"3871842e",
  1832 => x"09810680",
  1833 => x"f2388813",
  1834 => x"0851b0ee",
  1835 => x"2dba9704",
  1836 => x"80ccc808",
  1837 => x"51881308",
  1838 => x"52712dba",
  1839 => x"9704810b",
  1840 => x"8814082b",
  1841 => x"80ccb408",
  1842 => x"3280ccb4",
  1843 => x"0cb9eb04",
  1844 => x"881380f5",
  1845 => x"2d81058b",
  1846 => x"1480f52d",
  1847 => x"53547174",
  1848 => x"24833880",
  1849 => x"54738814",
  1850 => x"81b72daf",
  1851 => x"cb2dba97",
  1852 => x"04750880",
  1853 => x"2ea43875",
  1854 => x"0851aea0",
  1855 => x"2d80c290",
  1856 => x"08810652",
  1857 => x"71802e8c",
  1858 => x"3880ccc8",
  1859 => x"08518416",
  1860 => x"0852712d",
  1861 => x"88165675",
  1862 => x"d8388054",
  1863 => x"800b80c2",
  1864 => x"a40c738f",
  1865 => x"0680c2a0",
  1866 => x"0ca05273",
  1867 => x"80ccc808",
  1868 => x"2e098106",
  1869 => x"993880cc",
  1870 => x"c408ff05",
  1871 => x"74327009",
  1872 => x"81057072",
  1873 => x"079f2a91",
  1874 => x"71315151",
  1875 => x"53537151",
  1876 => x"82f82d81",
  1877 => x"14548e74",
  1878 => x"25c23880",
  1879 => x"c28c0852",
  1880 => x"7180c290",
  1881 => x"0c029805",
  1882 => x"0d040000",
  1883 => x"00ffffff",
  1884 => x"ff00ffff",
  1885 => x"ffff00ff",
  1886 => x"ffffff00",
  1887 => x"4f4b0000",
  1888 => x"52657365",
  1889 => x"74000000",
  1890 => x"53617665",
  1891 => x"20736574",
  1892 => x"74696e67",
  1893 => x"73000000",
  1894 => x"5363616e",
  1895 => x"6c696e65",
  1896 => x"73000000",
  1897 => x"41756469",
  1898 => x"6f20566f",
  1899 => x"6c756d65",
  1900 => x"00000000",
  1901 => x"4c6f6164",
  1902 => x"20524f4d",
  1903 => x"20100000",
  1904 => x"45786974",
  1905 => x"00000000",
  1906 => x"464d2064",
  1907 => x"69736162",
  1908 => x"6c650000",
  1909 => x"464d2065",
  1910 => x"6e61626c",
  1911 => x"65000000",
  1912 => x"50534720",
  1913 => x"64697361",
  1914 => x"626c6500",
  1915 => x"50534720",
  1916 => x"656e6162",
  1917 => x"6c650000",
  1918 => x"4a6f7973",
  1919 => x"7469636b",
  1920 => x"20737761",
  1921 => x"70000000",
  1922 => x"4a6f7973",
  1923 => x"7469636b",
  1924 => x"206e6f72",
  1925 => x"6d616c00",
  1926 => x"56474120",
  1927 => x"2d203331",
  1928 => x"4b487a00",
  1929 => x"5456202d",
  1930 => x"2031354b",
  1931 => x"487a0000",
  1932 => x"4261636b",
  1933 => x"00000000",
  1934 => x"4c6f6164",
  1935 => x"20457272",
  1936 => x"6f722100",
  1937 => x"46504741",
  1938 => x"47454e20",
  1939 => x"43464700",
  1940 => x"496e6974",
  1941 => x"69616c69",
  1942 => x"7a696e67",
  1943 => x"20534420",
  1944 => x"63617264",
  1945 => x"0a000000",
  1946 => x"424f4f54",
  1947 => x"20202020",
  1948 => x"47454e00",
  1949 => x"43617264",
  1950 => x"20696e69",
  1951 => x"74206661",
  1952 => x"696c6564",
  1953 => x"0a000000",
  1954 => x"4d425220",
  1955 => x"6661696c",
  1956 => x"0a000000",
  1957 => x"46415431",
  1958 => x"36202020",
  1959 => x"00000000",
  1960 => x"46415433",
  1961 => x"32202020",
  1962 => x"00000000",
  1963 => x"4e6f2070",
  1964 => x"61727469",
  1965 => x"74696f6e",
  1966 => x"20736967",
  1967 => x"0a000000",
  1968 => x"42616420",
  1969 => x"70617274",
  1970 => x"0a000000",
  1971 => x"53444843",
  1972 => x"20657272",
  1973 => x"6f72210a",
  1974 => x"00000000",
  1975 => x"53442069",
  1976 => x"6e69742e",
  1977 => x"2e2e0a00",
  1978 => x"53442063",
  1979 => x"61726420",
  1980 => x"72657365",
  1981 => x"74206661",
  1982 => x"696c6564",
  1983 => x"210a0000",
  1984 => x"57726974",
  1985 => x"65206661",
  1986 => x"696c6564",
  1987 => x"0a000000",
  1988 => x"52656164",
  1989 => x"20666169",
  1990 => x"6c65640a",
  1991 => x"00000000",
  1992 => x"16200000",
  1993 => x"14200000",
  1994 => x"15200000",
  1995 => x"00000002",
  1996 => x"00000000",
  1997 => x"00000002",
  1998 => x"00001d80",
  1999 => x"000004ff",
  2000 => x"00000002",
  2001 => x"00001d88",
  2002 => x"000003c4",
  2003 => x"00000003",
  2004 => x"00001fd0",
  2005 => x"00000002",
  2006 => x"00000001",
  2007 => x"00001d98",
  2008 => x"00000001",
  2009 => x"00000003",
  2010 => x"00001fc8",
  2011 => x"00000002",
  2012 => x"00000005",
  2013 => x"00001da4",
  2014 => x"00000007",
  2015 => x"00000003",
  2016 => x"00001fc0",
  2017 => x"00000002",
  2018 => x"00000003",
  2019 => x"00001fb8",
  2020 => x"00000002",
  2021 => x"00000002",
  2022 => x"00001db4",
  2023 => x"000007d3",
  2024 => x"00000002",
  2025 => x"00001dc0",
  2026 => x"00001787",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00001dc8",
  2031 => x"00001dd4",
  2032 => x"00001de0",
  2033 => x"00001dec",
  2034 => x"00001df8",
  2035 => x"00001e08",
  2036 => x"00001e18",
  2037 => x"00001e24",
  2038 => x"00000002",
  2039 => x"00002140",
  2040 => x"00000591",
  2041 => x"00000002",
  2042 => x"0000215e",
  2043 => x"00000591",
  2044 => x"00000002",
  2045 => x"0000217c",
  2046 => x"00000591",
  2047 => x"00000002",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

