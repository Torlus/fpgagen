-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM1 is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM1;

architecture arch of CtrlROM_ROM1 is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b80c1",
     9 => x"fc080b0b",
    10 => x"80c28008",
    11 => x"0b0b80c2",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c2840c0b",
    16 => x"0b80c280",
    17 => x"0c0b0b80",
    18 => x"c1fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbad8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c1fc70",
    57 => x"80ccb827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5190df",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c2",
    65 => x"8c0c9f0b",
    66 => x"80c2900c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c29008ff",
    70 => x"0580c290",
    71 => x"0c80c290",
    72 => x"088025e8",
    73 => x"3880c28c",
    74 => x"08ff0580",
    75 => x"c28c0c80",
    76 => x"c28c0880",
    77 => x"25d03802",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"80c28c08",
    97 => x"25913882",
    98 => x"bc2d80c2",
    99 => x"8c08ff05",
   100 => x"80c28c0c",
   101 => x"82fe0480",
   102 => x"c28c0880",
   103 => x"c2900853",
   104 => x"51728a2e",
   105 => x"098106be",
   106 => x"38715171",
   107 => x"9f24a438",
   108 => x"80c28c08",
   109 => x"a02911f8",
   110 => x"80115151",
   111 => x"a0713480",
   112 => x"c2900881",
   113 => x"0580c290",
   114 => x"0c80c290",
   115 => x"08519f71",
   116 => x"25de3880",
   117 => x"0b80c290",
   118 => x"0c80c28c",
   119 => x"08810580",
   120 => x"c28c0c83",
   121 => x"fc0470a0",
   122 => x"2912f880",
   123 => x"11515172",
   124 => x"713480c2",
   125 => x"90088105",
   126 => x"80c2900c",
   127 => x"80c29008",
   128 => x"a02e0981",
   129 => x"06913880",
   130 => x"0b80c290",
   131 => x"0c80c28c",
   132 => x"08810580",
   133 => x"c28c0c02",
   134 => x"8c050d04",
   135 => x"02e8050d",
   136 => x"77795656",
   137 => x"880bfc16",
   138 => x"77712c8f",
   139 => x"06545254",
   140 => x"80537272",
   141 => x"25953871",
   142 => x"53fbe014",
   143 => x"51877134",
   144 => x"8114ff14",
   145 => x"545472f1",
   146 => x"387153f9",
   147 => x"1576712c",
   148 => x"87065351",
   149 => x"71802e8b",
   150 => x"38fbe014",
   151 => x"51717134",
   152 => x"81145472",
   153 => x"8e249538",
   154 => x"8f733153",
   155 => x"fbe01451",
   156 => x"a0713481",
   157 => x"14ff1454",
   158 => x"5472f138",
   159 => x"0298050d",
   160 => x"0402ec05",
   161 => x"0d800b80",
   162 => x"c2940cf6",
   163 => x"8c08f690",
   164 => x"0871882c",
   165 => x"565481ff",
   166 => x"06527372",
   167 => x"25893871",
   168 => x"54820b80",
   169 => x"c2940c72",
   170 => x"882c7381",
   171 => x"ff065455",
   172 => x"7473258d",
   173 => x"387280c2",
   174 => x"94088407",
   175 => x"80c2940c",
   176 => x"5573842b",
   177 => x"87e87125",
   178 => x"83713170",
   179 => x"0b0b0bbe",
   180 => x"980c8171",
   181 => x"2bf6880c",
   182 => x"fea413ff",
   183 => x"122c7888",
   184 => x"29ff9405",
   185 => x"70812c80",
   186 => x"c2940852",
   187 => x"58525551",
   188 => x"52547680",
   189 => x"2e853870",
   190 => x"81075170",
   191 => x"f6940c71",
   192 => x"098105f6",
   193 => x"800c7209",
   194 => x"8105f684",
   195 => x"0c029405",
   196 => x"0d0402f4",
   197 => x"050d7453",
   198 => x"72708105",
   199 => x"5480f52d",
   200 => x"5271802e",
   201 => x"89387151",
   202 => x"82f82d86",
   203 => x"9804028c",
   204 => x"050d0402",
   205 => x"f4050d74",
   206 => x"70820680",
   207 => x"cc9c0cbe",
   208 => x"b8718106",
   209 => x"53535370",
   210 => x"881381b7",
   211 => x"2d981273",
   212 => x"822a7081",
   213 => x"06515252",
   214 => x"70881381",
   215 => x"b72d9812",
   216 => x"73832a70",
   217 => x"81065152",
   218 => x"52708813",
   219 => x"81b72d72",
   220 => x"842a7081",
   221 => x"06515372",
   222 => x"941381b7",
   223 => x"2d7080c1",
   224 => x"fc0c028c",
   225 => x"050d0402",
   226 => x"f8050dbc",
   227 => x"b05280c2",
   228 => x"98519ed4",
   229 => x"2d80c1fc",
   230 => x"08802ea3",
   231 => x"3880c5b0",
   232 => x"5280c298",
   233 => x"51a1a12d",
   234 => x"80c5b008",
   235 => x"80c2a40c",
   236 => x"80c5b008",
   237 => x"fec00c80",
   238 => x"c5b00851",
   239 => x"86b32d02",
   240 => x"88050d04",
   241 => x"02f0050d",
   242 => x"80519488",
   243 => x"2dbcb052",
   244 => x"80c29851",
   245 => x"9ed42d80",
   246 => x"c1fc0880",
   247 => x"2eaa3880",
   248 => x"c2a40880",
   249 => x"c5b00c80",
   250 => x"c5b45480",
   251 => x"fd538074",
   252 => x"70840556",
   253 => x"0cff1353",
   254 => x"728025f2",
   255 => x"3880c5b0",
   256 => x"5280c298",
   257 => x"51a1ca2d",
   258 => x"0290050d",
   259 => x"0402d805",
   260 => x"0d800bbe",
   261 => x"9c0c80c2",
   262 => x"a408fec0",
   263 => x"0c810bfe",
   264 => x"c40c840b",
   265 => x"fec40c7b",
   266 => x"5280c298",
   267 => x"519ed42d",
   268 => x"80c1fc08",
   269 => x"5380c1fc",
   270 => x"08802e81",
   271 => x"b83880c2",
   272 => x"9c085580",
   273 => x"0bff1657",
   274 => x"5975792e",
   275 => x"8b388119",
   276 => x"76812a57",
   277 => x"5975f738",
   278 => x"f7195974",
   279 => x"b080802e",
   280 => x"09810689",
   281 => x"38820bfe",
   282 => x"dc0c8984",
   283 => x"04749880",
   284 => x"802e0981",
   285 => x"06893881",
   286 => x"0bfedc0c",
   287 => x"89840480",
   288 => x"0bfedc0c",
   289 => x"815a8075",
   290 => x"2580e338",
   291 => x"78527551",
   292 => x"849c2d80",
   293 => x"c5b05280",
   294 => x"c29851a1",
   295 => x"a12d80c1",
   296 => x"fc08802e",
   297 => x"a83880c5",
   298 => x"b05883fc",
   299 => x"57777084",
   300 => x"05590870",
   301 => x"83ffff06",
   302 => x"71902afe",
   303 => x"c80cfec8",
   304 => x"0cfc1858",
   305 => x"53768025",
   306 => x"e43889d5",
   307 => x"0480c1fc",
   308 => x"085a8480",
   309 => x"5580c298",
   310 => x"51a0f12d",
   311 => x"fc801581",
   312 => x"17575574",
   313 => x"8024ffa4",
   314 => x"3879802e",
   315 => x"8638820b",
   316 => x"be9c0c79",
   317 => x"537280c1",
   318 => x"fc0c02a8",
   319 => x"050d0402",
   320 => x"fc050dae",
   321 => x"f52dfec4",
   322 => x"5181710c",
   323 => x"82710c02",
   324 => x"84050d04",
   325 => x"02f4050d",
   326 => x"74767853",
   327 => x"54528071",
   328 => x"25973872",
   329 => x"70810554",
   330 => x"80f52d72",
   331 => x"70810554",
   332 => x"81b72dff",
   333 => x"115170eb",
   334 => x"38807281",
   335 => x"b72d028c",
   336 => x"050d0402",
   337 => x"e8050d77",
   338 => x"56807056",
   339 => x"54737624",
   340 => x"b63880cb",
   341 => x"c008742e",
   342 => x"ae387351",
   343 => x"9c992d80",
   344 => x"c1fc0880",
   345 => x"c1fc0809",
   346 => x"81057080",
   347 => x"c1fc0807",
   348 => x"9f2a7705",
   349 => x"81175757",
   350 => x"53537476",
   351 => x"24893880",
   352 => x"cbc00874",
   353 => x"26d43872",
   354 => x"80c1fc0c",
   355 => x"0298050d",
   356 => x"0402f405",
   357 => x"0d80c0f8",
   358 => x"0815518a",
   359 => x"c32d80c1",
   360 => x"fc08802e",
   361 => x"ac388b53",
   362 => x"80c1fc08",
   363 => x"5280c9b0",
   364 => x"518a942d",
   365 => x"80c9b051",
   366 => x"888d2d80",
   367 => x"c1fc0880",
   368 => x"2e8f38be",
   369 => x"a051b0dc",
   370 => x"2daef52d",
   371 => x"80518bdd",
   372 => x"0480c0fc",
   373 => x"51b0dc2d",
   374 => x"aee12d81",
   375 => x"5185812d",
   376 => x"028c050d",
   377 => x"0402dc05",
   378 => x"0d80705a",
   379 => x"557480c0",
   380 => x"f80825b4",
   381 => x"3880cbc0",
   382 => x"08752eac",
   383 => x"3878519c",
   384 => x"992d80c1",
   385 => x"fc080981",
   386 => x"057080c1",
   387 => x"fc08079f",
   388 => x"2a760581",
   389 => x"1b5b5654",
   390 => x"7480c0f8",
   391 => x"08258938",
   392 => x"80cbc008",
   393 => x"7926d638",
   394 => x"80557880",
   395 => x"cbc00827",
   396 => x"81d93878",
   397 => x"519c992d",
   398 => x"80c1fc08",
   399 => x"802e81ab",
   400 => x"3880c1fc",
   401 => x"088b0580",
   402 => x"f52d7084",
   403 => x"2a708106",
   404 => x"77107884",
   405 => x"2b80c9b0",
   406 => x"0b80f52d",
   407 => x"5c5c5351",
   408 => x"55567380",
   409 => x"2e80ca38",
   410 => x"7416822b",
   411 => x"8eaf0bbf",
   412 => x"cc120c54",
   413 => x"77753110",
   414 => x"80c2a811",
   415 => x"55569074",
   416 => x"70810556",
   417 => x"81b72da0",
   418 => x"7481b72d",
   419 => x"7681ff06",
   420 => x"81165854",
   421 => x"73802e8a",
   422 => x"389c5380",
   423 => x"c9b0528d",
   424 => x"a9048b53",
   425 => x"80c1fc08",
   426 => x"5280c2aa",
   427 => x"16518de3",
   428 => x"04741682",
   429 => x"2b8b910b",
   430 => x"bfcc120c",
   431 => x"547681ff",
   432 => x"06811658",
   433 => x"5473802e",
   434 => x"8a389c53",
   435 => x"80c9b052",
   436 => x"8dda048b",
   437 => x"5380c1fc",
   438 => x"08527775",
   439 => x"311080c2",
   440 => x"a8055176",
   441 => x"558a942d",
   442 => x"8e800474",
   443 => x"90297531",
   444 => x"701080c2",
   445 => x"a8055154",
   446 => x"80c1fc08",
   447 => x"7481b72d",
   448 => x"81195974",
   449 => x"8b24a338",
   450 => x"8caa0474",
   451 => x"90297531",
   452 => x"701080c2",
   453 => x"a8058c77",
   454 => x"31575154",
   455 => x"807481b7",
   456 => x"2d9e14ff",
   457 => x"16565474",
   458 => x"f33802a4",
   459 => x"050d0402",
   460 => x"fc050d80",
   461 => x"c0f80813",
   462 => x"518ac32d",
   463 => x"80c1fc08",
   464 => x"802e8938",
   465 => x"80c1fc08",
   466 => x"5194882d",
   467 => x"800b80c0",
   468 => x"f80c8be5",
   469 => x"2dafb92d",
   470 => x"0284050d",
   471 => x"0402fc05",
   472 => x"0d725170",
   473 => x"fd2eb038",
   474 => x"70fd248a",
   475 => x"3870fc2e",
   476 => x"80cc388f",
   477 => x"c80470fe",
   478 => x"2eb73870",
   479 => x"ff2e0981",
   480 => x"0680c538",
   481 => x"80c0f808",
   482 => x"5170802e",
   483 => x"bb38ff11",
   484 => x"80c0f80c",
   485 => x"8fc80480",
   486 => x"c0f808f0",
   487 => x"057080c0",
   488 => x"f80c5170",
   489 => x"8025a138",
   490 => x"800b80c0",
   491 => x"f80c8fc8",
   492 => x"0480c0f8",
   493 => x"08810580",
   494 => x"c0f80c8f",
   495 => x"c80480c0",
   496 => x"f8089005",
   497 => x"80c0f80c",
   498 => x"8be52daf",
   499 => x"b92d0284",
   500 => x"050d0402",
   501 => x"fc050d80",
   502 => x"0b80c0f8",
   503 => x"0c8be52d",
   504 => x"bfc451b0",
   505 => x"dc2d0284",
   506 => x"050d04be",
   507 => x"e40b80f5",
   508 => x"2d80c1fc",
   509 => x"0c0402fc",
   510 => x"050d7287",
   511 => x"065170be",
   512 => x"e40b81b7",
   513 => x"2d028405",
   514 => x"0d0402f8",
   515 => x"050d80cc",
   516 => x"9c088206",
   517 => x"bec00b80",
   518 => x"f52d5252",
   519 => x"70802e85",
   520 => x"38718107",
   521 => x"52bed80b",
   522 => x"80f52d51",
   523 => x"70802e85",
   524 => x"38718407",
   525 => x"52bef00b",
   526 => x"80f52d51",
   527 => x"70802e85",
   528 => x"38718807",
   529 => x"52befc0b",
   530 => x"80f52d51",
   531 => x"70802e85",
   532 => x"38719007",
   533 => x"527180c1",
   534 => x"fc0c0288",
   535 => x"050d0402",
   536 => x"f0050d80",
   537 => x"0bbe9c0c",
   538 => x"87538051",
   539 => x"86b32d72",
   540 => x"518ff62d",
   541 => x"810bfec4",
   542 => x"0c840bfe",
   543 => x"c40c830b",
   544 => x"fecc0cbc",
   545 => x"bc518692",
   546 => x"2d8452a6",
   547 => x"902d95ae",
   548 => x"2d80c1fc",
   549 => x"08802e86",
   550 => x"38fe5291",
   551 => x"a604ff12",
   552 => x"52718024",
   553 => x"e6387180",
   554 => x"2e828d38",
   555 => x"acae2dae",
   556 => x"d52dac91",
   557 => x"2dac912d",
   558 => x"81f92d81",
   559 => x"5185812d",
   560 => x"ac912dac",
   561 => x"912d8151",
   562 => x"85812d87",
   563 => x"872dbcd4",
   564 => x"51888d2d",
   565 => x"80c1fc08",
   566 => x"802e9438",
   567 => x"bea051b0",
   568 => x"dc2d8051",
   569 => x"85812d82",
   570 => x"0bbe9c0c",
   571 => x"91fa0480",
   572 => x"c1fc0851",
   573 => x"8fd32dae",
   574 => x"e12dacc7",
   575 => x"2db0ef2d",
   576 => x"80c1fc08",
   577 => x"80cca008",
   578 => x"882b80cc",
   579 => x"a40807fe",
   580 => x"d80c5490",
   581 => x"8a2d80c1",
   582 => x"fc0880c2",
   583 => x"a4082ea5",
   584 => x"3880c1fc",
   585 => x"0880c2a4",
   586 => x"0c80c1fc",
   587 => x"08fec00c",
   588 => x"84527351",
   589 => x"85812dac",
   590 => x"912dac91",
   591 => x"2dff1252",
   592 => x"718025ee",
   593 => x"388551ae",
   594 => x"8e2d80c1",
   595 => x"fc08812a",
   596 => x"70810651",
   597 => x"5271802e",
   598 => x"9538ff13",
   599 => x"7009709f",
   600 => x"2c720670",
   601 => x"54525353",
   602 => x"8ff62daf",
   603 => x"b92d8651",
   604 => x"ae8e2d80",
   605 => x"c1fc0881",
   606 => x"2a708106",
   607 => x"51527180",
   608 => x"2e933881",
   609 => x"13538773",
   610 => x"25833887",
   611 => x"5372518f",
   612 => x"f62dafb9",
   613 => x"2d8feb2d",
   614 => x"80c1fc08",
   615 => x"fed40c73",
   616 => x"802e8c38",
   617 => x"be9c0888",
   618 => x"07fec40c",
   619 => x"91fa04be",
   620 => x"9c08fec4",
   621 => x"0c91fa04",
   622 => x"bce05186",
   623 => x"922d800b",
   624 => x"80c1fc0c",
   625 => x"0290050d",
   626 => x"0402e805",
   627 => x"0d77797b",
   628 => x"58555580",
   629 => x"53727625",
   630 => x"a3387470",
   631 => x"81055680",
   632 => x"f52d7470",
   633 => x"81055680",
   634 => x"f52d5252",
   635 => x"71712e86",
   636 => x"38815193",
   637 => x"fe048113",
   638 => x"5393d504",
   639 => x"80517080",
   640 => x"c1fc0c02",
   641 => x"98050d04",
   642 => x"02ec050d",
   643 => x"76557480",
   644 => x"2e80c238",
   645 => x"9a1580e0",
   646 => x"2d51aad4",
   647 => x"2d80c1fc",
   648 => x"0880c1fc",
   649 => x"0880cbe0",
   650 => x"0c80c1fc",
   651 => x"08545480",
   652 => x"cbbc0880",
   653 => x"2e9a3894",
   654 => x"1580e02d",
   655 => x"51aad42d",
   656 => x"80c1fc08",
   657 => x"902b83ff",
   658 => x"f00a0670",
   659 => x"75075153",
   660 => x"7280cbe0",
   661 => x"0c80cbe0",
   662 => x"08537280",
   663 => x"2e9d3880",
   664 => x"cbb408fe",
   665 => x"14712980",
   666 => x"cbc80805",
   667 => x"80cbe40c",
   668 => x"70842b80",
   669 => x"cbc00c54",
   670 => x"95a90480",
   671 => x"cbcc0880",
   672 => x"cbe00c80",
   673 => x"cbd00880",
   674 => x"cbe40c80",
   675 => x"cbbc0880",
   676 => x"2e8b3880",
   677 => x"cbb40884",
   678 => x"2b5395a4",
   679 => x"0480cbd4",
   680 => x"08842b53",
   681 => x"7280cbc0",
   682 => x"0c029405",
   683 => x"0d0402d8",
   684 => x"050d800b",
   685 => x"80cbbc0c",
   686 => x"80c5b052",
   687 => x"8051a980",
   688 => x"2d80c1fc",
   689 => x"085480c1",
   690 => x"fc088c38",
   691 => x"bcf45186",
   692 => x"922d7355",
   693 => x"9b960480",
   694 => x"56810b80",
   695 => x"cbe80c88",
   696 => x"53bd8052",
   697 => x"80c5e651",
   698 => x"93c92d80",
   699 => x"c1fc0876",
   700 => x"2e098106",
   701 => x"893880c1",
   702 => x"fc0880cb",
   703 => x"e80c8853",
   704 => x"bd8c5280",
   705 => x"c6825193",
   706 => x"c92d80c1",
   707 => x"fc088938",
   708 => x"80c1fc08",
   709 => x"80cbe80c",
   710 => x"80cbe808",
   711 => x"802e8180",
   712 => x"3880c8f6",
   713 => x"0b80f52d",
   714 => x"80c8f70b",
   715 => x"80f52d71",
   716 => x"982b7190",
   717 => x"2b0780c8",
   718 => x"f80b80f5",
   719 => x"2d70882b",
   720 => x"720780c8",
   721 => x"f90b80f5",
   722 => x"2d710780",
   723 => x"c9ae0b80",
   724 => x"f52d80c9",
   725 => x"af0b80f5",
   726 => x"2d71882b",
   727 => x"07535f54",
   728 => x"525a5657",
   729 => x"557381ab",
   730 => x"aa2e0981",
   731 => x"068e3875",
   732 => x"51aaa32d",
   733 => x"80c1fc08",
   734 => x"56978904",
   735 => x"7382d4d5",
   736 => x"2e8738bd",
   737 => x"985197d2",
   738 => x"0480c5b0",
   739 => x"527551a9",
   740 => x"802d80c1",
   741 => x"fc085580",
   742 => x"c1fc0880",
   743 => x"2e83f738",
   744 => x"8853bd8c",
   745 => x"5280c682",
   746 => x"5193c92d",
   747 => x"80c1fc08",
   748 => x"8a38810b",
   749 => x"80cbbc0c",
   750 => x"97d80488",
   751 => x"53bd8052",
   752 => x"80c5e651",
   753 => x"93c92d80",
   754 => x"c1fc0880",
   755 => x"2e8a38bd",
   756 => x"ac518692",
   757 => x"2d98b704",
   758 => x"80c9ae0b",
   759 => x"80f52d54",
   760 => x"7380d52e",
   761 => x"09810680",
   762 => x"ce3880c9",
   763 => x"af0b80f5",
   764 => x"2d547381",
   765 => x"aa2e0981",
   766 => x"06bd3880",
   767 => x"0b80c5b0",
   768 => x"0b80f52d",
   769 => x"56547481",
   770 => x"e92e8338",
   771 => x"81547481",
   772 => x"eb2e8c38",
   773 => x"80557375",
   774 => x"2e098106",
   775 => x"82f83880",
   776 => x"c5bb0b80",
   777 => x"f52d5574",
   778 => x"8e3880c5",
   779 => x"bc0b80f5",
   780 => x"2d547382",
   781 => x"2e863880",
   782 => x"559b9604",
   783 => x"80c5bd0b",
   784 => x"80f52d70",
   785 => x"80cbb40c",
   786 => x"ff0580cb",
   787 => x"b80c80c5",
   788 => x"be0b80f5",
   789 => x"2d80c5bf",
   790 => x"0b80f52d",
   791 => x"58760577",
   792 => x"82802905",
   793 => x"7080cbc4",
   794 => x"0c80c5c0",
   795 => x"0b80f52d",
   796 => x"7080cbd8",
   797 => x"0c80cbbc",
   798 => x"08595758",
   799 => x"76802e81",
   800 => x"b6388853",
   801 => x"bd8c5280",
   802 => x"c6825193",
   803 => x"c92d80c1",
   804 => x"fc088282",
   805 => x"3880cbb4",
   806 => x"0870842b",
   807 => x"80cbc00c",
   808 => x"7080cbd4",
   809 => x"0c80c5d5",
   810 => x"0b80f52d",
   811 => x"80c5d40b",
   812 => x"80f52d71",
   813 => x"82802905",
   814 => x"80c5d60b",
   815 => x"80f52d70",
   816 => x"84808029",
   817 => x"1280c5d7",
   818 => x"0b80f52d",
   819 => x"7081800a",
   820 => x"29127080",
   821 => x"cbdc0c80",
   822 => x"cbd80871",
   823 => x"2980cbc4",
   824 => x"08057080",
   825 => x"cbc80c80",
   826 => x"c5dd0b80",
   827 => x"f52d80c5",
   828 => x"dc0b80f5",
   829 => x"2d718280",
   830 => x"290580c5",
   831 => x"de0b80f5",
   832 => x"2d708480",
   833 => x"80291280",
   834 => x"c5df0b80",
   835 => x"f52d7098",
   836 => x"2b81f00a",
   837 => x"06720570",
   838 => x"80cbcc0c",
   839 => x"fe117e29",
   840 => x"770580cb",
   841 => x"d00c5259",
   842 => x"5243545e",
   843 => x"51525952",
   844 => x"5d575957",
   845 => x"9b8f0480",
   846 => x"c5c20b80",
   847 => x"f52d80c5",
   848 => x"c10b80f5",
   849 => x"2d718280",
   850 => x"29057080",
   851 => x"cbc00c70",
   852 => x"a02983ff",
   853 => x"0570892a",
   854 => x"7080cbd4",
   855 => x"0c80c5c7",
   856 => x"0b80f52d",
   857 => x"80c5c60b",
   858 => x"80f52d71",
   859 => x"82802905",
   860 => x"7080cbdc",
   861 => x"0c7b7129",
   862 => x"1e7080cb",
   863 => x"d00c7d80",
   864 => x"cbcc0c73",
   865 => x"0580cbc8",
   866 => x"0c555e51",
   867 => x"51555580",
   868 => x"5194882d",
   869 => x"81557480",
   870 => x"c1fc0c02",
   871 => x"a8050d04",
   872 => x"02ec050d",
   873 => x"7670872c",
   874 => x"7180ff06",
   875 => x"55565480",
   876 => x"cbbc088a",
   877 => x"3873882c",
   878 => x"7481ff06",
   879 => x"545580c5",
   880 => x"b05280cb",
   881 => x"c4081551",
   882 => x"a9802d80",
   883 => x"c1fc0854",
   884 => x"80c1fc08",
   885 => x"802eb838",
   886 => x"80cbbc08",
   887 => x"802e9a38",
   888 => x"72842980",
   889 => x"c5b00570",
   890 => x"085253aa",
   891 => x"a32d80c1",
   892 => x"fc08f00a",
   893 => x"06539c8d",
   894 => x"04721080",
   895 => x"c5b00570",
   896 => x"80e02d52",
   897 => x"53aad42d",
   898 => x"80c1fc08",
   899 => x"53725473",
   900 => x"80c1fc0c",
   901 => x"0294050d",
   902 => x"0402e005",
   903 => x"0d797084",
   904 => x"2c80cbe4",
   905 => x"0805718f",
   906 => x"06525553",
   907 => x"728a3880",
   908 => x"c5b05273",
   909 => x"51a9802d",
   910 => x"72a02980",
   911 => x"c5b00554",
   912 => x"807480f5",
   913 => x"2d565374",
   914 => x"732e8338",
   915 => x"81537481",
   916 => x"e52e81f4",
   917 => x"38817074",
   918 => x"06545872",
   919 => x"802e81e8",
   920 => x"388b1480",
   921 => x"f52d7083",
   922 => x"2a790658",
   923 => x"56769b38",
   924 => x"80c1ac08",
   925 => x"53728938",
   926 => x"7280c9b0",
   927 => x"0b81b72d",
   928 => x"7680c1ac",
   929 => x"0c73539e",
   930 => x"ca04758f",
   931 => x"2e098106",
   932 => x"81b63874",
   933 => x"9f068d29",
   934 => x"80c9a311",
   935 => x"51538114",
   936 => x"80f52d73",
   937 => x"70810555",
   938 => x"81b72d83",
   939 => x"1480f52d",
   940 => x"73708105",
   941 => x"5581b72d",
   942 => x"851480f5",
   943 => x"2d737081",
   944 => x"055581b7",
   945 => x"2d871480",
   946 => x"f52d7370",
   947 => x"81055581",
   948 => x"b72d8914",
   949 => x"80f52d73",
   950 => x"70810555",
   951 => x"81b72d8e",
   952 => x"1480f52d",
   953 => x"73708105",
   954 => x"5581b72d",
   955 => x"901480f5",
   956 => x"2d737081",
   957 => x"055581b7",
   958 => x"2d921480",
   959 => x"f52d7370",
   960 => x"81055581",
   961 => x"b72d9414",
   962 => x"80f52d73",
   963 => x"70810555",
   964 => x"81b72d96",
   965 => x"1480f52d",
   966 => x"73708105",
   967 => x"5581b72d",
   968 => x"981480f5",
   969 => x"2d737081",
   970 => x"055581b7",
   971 => x"2d9c1480",
   972 => x"f52d7370",
   973 => x"81055581",
   974 => x"b72d9e14",
   975 => x"80f52d73",
   976 => x"81b72d77",
   977 => x"80c1ac0c",
   978 => x"80537280",
   979 => x"c1fc0c02",
   980 => x"a0050d04",
   981 => x"02cc050d",
   982 => x"7e605e5a",
   983 => x"800b80cb",
   984 => x"e00880cb",
   985 => x"e408595c",
   986 => x"56805880",
   987 => x"cbc00878",
   988 => x"2e81b838",
   989 => x"778f06a0",
   990 => x"17575473",
   991 => x"913880c5",
   992 => x"b0527651",
   993 => x"811757a9",
   994 => x"802d80c5",
   995 => x"b0568076",
   996 => x"80f52d56",
   997 => x"5474742e",
   998 => x"83388154",
   999 => x"7481e52e",
  1000 => x"80fd3881",
  1001 => x"70750655",
  1002 => x"5c73802e",
  1003 => x"80f1388b",
  1004 => x"1680f52d",
  1005 => x"98065978",
  1006 => x"80e5388b",
  1007 => x"537c5275",
  1008 => x"5193c92d",
  1009 => x"80c1fc08",
  1010 => x"80d5389c",
  1011 => x"160851aa",
  1012 => x"a32d80c1",
  1013 => x"fc08841b",
  1014 => x"0c9a1680",
  1015 => x"e02d51aa",
  1016 => x"d42d80c1",
  1017 => x"fc0880c1",
  1018 => x"fc08881c",
  1019 => x"0c80c1fc",
  1020 => x"08555580",
  1021 => x"cbbc0880",
  1022 => x"2e993894",
  1023 => x"1680e02d",
  1024 => x"51aad42d",
  1025 => x"80c1fc08",
  1026 => x"902b83ff",
  1027 => x"f00a0670",
  1028 => x"16515473",
  1029 => x"881b0c78",
  1030 => x"7a0c7b54",
  1031 => x"a0e70481",
  1032 => x"185880cb",
  1033 => x"c0087826",
  1034 => x"feca3880",
  1035 => x"cbbc0880",
  1036 => x"2eb3387a",
  1037 => x"519ba02d",
  1038 => x"80c1fc08",
  1039 => x"80c1fc08",
  1040 => x"80ffffff",
  1041 => x"f806555b",
  1042 => x"7380ffff",
  1043 => x"fff82e95",
  1044 => x"3880c1fc",
  1045 => x"08fe0580",
  1046 => x"cbb40829",
  1047 => x"80cbc808",
  1048 => x"05579ee9",
  1049 => x"04805473",
  1050 => x"80c1fc0c",
  1051 => x"02b4050d",
  1052 => x"0402f405",
  1053 => x"0d747008",
  1054 => x"8105710c",
  1055 => x"700880cb",
  1056 => x"b8080653",
  1057 => x"53718f38",
  1058 => x"88130851",
  1059 => x"9ba02d80",
  1060 => x"c1fc0888",
  1061 => x"140c810b",
  1062 => x"80c1fc0c",
  1063 => x"028c050d",
  1064 => x"0402f005",
  1065 => x"0d758811",
  1066 => x"08fe0580",
  1067 => x"cbb40829",
  1068 => x"80cbc808",
  1069 => x"11720880",
  1070 => x"cbb80806",
  1071 => x"05795553",
  1072 => x"5454a980",
  1073 => x"2d029005",
  1074 => x"0d0402f0",
  1075 => x"050d7588",
  1076 => x"1108fe05",
  1077 => x"80cbb408",
  1078 => x"2980cbc8",
  1079 => x"08117208",
  1080 => x"80cbb808",
  1081 => x"06057955",
  1082 => x"535454a7",
  1083 => x"be2d0290",
  1084 => x"050d0402",
  1085 => x"f4050dd4",
  1086 => x"5281ff72",
  1087 => x"0c710853",
  1088 => x"81ff720c",
  1089 => x"72882b83",
  1090 => x"fe800672",
  1091 => x"087081ff",
  1092 => x"06515253",
  1093 => x"81ff720c",
  1094 => x"72710788",
  1095 => x"2b720870",
  1096 => x"81ff0651",
  1097 => x"525381ff",
  1098 => x"720c7271",
  1099 => x"07882b72",
  1100 => x"087081ff",
  1101 => x"06720780",
  1102 => x"c1fc0c52",
  1103 => x"53028c05",
  1104 => x"0d0402f4",
  1105 => x"050d7476",
  1106 => x"7181ff06",
  1107 => x"d40c5353",
  1108 => x"80cbec08",
  1109 => x"85387189",
  1110 => x"2b527198",
  1111 => x"2ad40c71",
  1112 => x"902a7081",
  1113 => x"ff06d40c",
  1114 => x"5171882a",
  1115 => x"7081ff06",
  1116 => x"d40c5171",
  1117 => x"81ff06d4",
  1118 => x"0c72902a",
  1119 => x"7081ff06",
  1120 => x"d40c51d4",
  1121 => x"087081ff",
  1122 => x"06515182",
  1123 => x"b8bf5270",
  1124 => x"81ff2e09",
  1125 => x"81069438",
  1126 => x"81ff0bd4",
  1127 => x"0cd40870",
  1128 => x"81ff06ff",
  1129 => x"14545151",
  1130 => x"71e53870",
  1131 => x"80c1fc0c",
  1132 => x"028c050d",
  1133 => x"0402fc05",
  1134 => x"0d81c751",
  1135 => x"81ff0bd4",
  1136 => x"0cff1151",
  1137 => x"708025f4",
  1138 => x"38028405",
  1139 => x"0d0402f0",
  1140 => x"050da3b5",
  1141 => x"2d8fcf53",
  1142 => x"805287fc",
  1143 => x"80f751a2",
  1144 => x"c22d80c1",
  1145 => x"fc085480",
  1146 => x"c1fc0881",
  1147 => x"2e098106",
  1148 => x"a43881ff",
  1149 => x"0bd40c82",
  1150 => x"0a52849c",
  1151 => x"80e951a2",
  1152 => x"c22d80c1",
  1153 => x"fc088b38",
  1154 => x"81ff0bd4",
  1155 => x"0c7353a4",
  1156 => x"9c04a3b5",
  1157 => x"2dff1353",
  1158 => x"72ffbd38",
  1159 => x"7280c1fc",
  1160 => x"0c029005",
  1161 => x"0d0402f4",
  1162 => x"050d81ff",
  1163 => x"0bd40c93",
  1164 => x"53805287",
  1165 => x"fc80c151",
  1166 => x"a2c22d80",
  1167 => x"c1fc088b",
  1168 => x"3881ff0b",
  1169 => x"d40c8153",
  1170 => x"a4d404a3",
  1171 => x"b52dff13",
  1172 => x"5372de38",
  1173 => x"7280c1fc",
  1174 => x"0c028c05",
  1175 => x"0d0402f0",
  1176 => x"050da3b5",
  1177 => x"2d83aa52",
  1178 => x"849c80c8",
  1179 => x"51a2c22d",
  1180 => x"80c1fc08",
  1181 => x"812e0981",
  1182 => x"069338a1",
  1183 => x"f32d80c1",
  1184 => x"fc0883ff",
  1185 => x"ff065372",
  1186 => x"83aa2e97",
  1187 => x"38a4a62d",
  1188 => x"a59e0481",
  1189 => x"54a68604",
  1190 => x"bdb85186",
  1191 => x"922d8054",
  1192 => x"a6860481",
  1193 => x"ff0bd40c",
  1194 => x"b153a3ce",
  1195 => x"2d80c1fc",
  1196 => x"08802e80",
  1197 => x"c2388052",
  1198 => x"87fc80fa",
  1199 => x"51a2c22d",
  1200 => x"80c1fc08",
  1201 => x"b23881ff",
  1202 => x"0bd40cd4",
  1203 => x"085381ff",
  1204 => x"0bd40c81",
  1205 => x"ff0bd40c",
  1206 => x"81ff0bd4",
  1207 => x"0c81ff0b",
  1208 => x"d40c7286",
  1209 => x"2a708106",
  1210 => x"80c1fc08",
  1211 => x"56515372",
  1212 => x"802e9338",
  1213 => x"a5930472",
  1214 => x"822eff9c",
  1215 => x"38ff1353",
  1216 => x"72ffa738",
  1217 => x"72547380",
  1218 => x"c1fc0c02",
  1219 => x"90050d04",
  1220 => x"02f0050d",
  1221 => x"810b80cb",
  1222 => x"ec0c8454",
  1223 => x"d008708f",
  1224 => x"2a708106",
  1225 => x"51515372",
  1226 => x"f33872d0",
  1227 => x"0ca3b52d",
  1228 => x"bdc85186",
  1229 => x"922dd008",
  1230 => x"708f2a70",
  1231 => x"81065151",
  1232 => x"5372f338",
  1233 => x"810bd00c",
  1234 => x"b1538052",
  1235 => x"84d480c0",
  1236 => x"51a2c22d",
  1237 => x"80c1fc08",
  1238 => x"812ea138",
  1239 => x"72822e09",
  1240 => x"81068c38",
  1241 => x"bdd45186",
  1242 => x"922d8053",
  1243 => x"a7b404ff",
  1244 => x"135372d6",
  1245 => x"38ff1454",
  1246 => x"73ffa138",
  1247 => x"a4de2d80",
  1248 => x"c1fc0880",
  1249 => x"cbec0c80",
  1250 => x"c1fc088b",
  1251 => x"38815287",
  1252 => x"fc80d051",
  1253 => x"a2c22d81",
  1254 => x"ff0bd40c",
  1255 => x"d008708f",
  1256 => x"2a708106",
  1257 => x"51515372",
  1258 => x"f33872d0",
  1259 => x"0c81ff0b",
  1260 => x"d40c8153",
  1261 => x"7280c1fc",
  1262 => x"0c029005",
  1263 => x"0d0402e8",
  1264 => x"050d7856",
  1265 => x"81ff0bd4",
  1266 => x"0cd00870",
  1267 => x"8f2a7081",
  1268 => x"06515153",
  1269 => x"72f33882",
  1270 => x"810bd00c",
  1271 => x"81ff0bd4",
  1272 => x"0c775287",
  1273 => x"fc80d851",
  1274 => x"a2c22d80",
  1275 => x"c1fc0880",
  1276 => x"2e8c38bd",
  1277 => x"ec518692",
  1278 => x"2d8153a8",
  1279 => x"f60481ff",
  1280 => x"0bd40c81",
  1281 => x"fe0bd40c",
  1282 => x"80ff5575",
  1283 => x"70840557",
  1284 => x"0870982a",
  1285 => x"d40c7090",
  1286 => x"2c7081ff",
  1287 => x"06d40c54",
  1288 => x"70882c70",
  1289 => x"81ff06d4",
  1290 => x"0c547081",
  1291 => x"ff06d40c",
  1292 => x"54ff1555",
  1293 => x"748025d3",
  1294 => x"3881ff0b",
  1295 => x"d40c81ff",
  1296 => x"0bd40c81",
  1297 => x"ff0bd40c",
  1298 => x"868da054",
  1299 => x"81ff0bd4",
  1300 => x"0cd40881",
  1301 => x"ff065574",
  1302 => x"8738ff14",
  1303 => x"5473ed38",
  1304 => x"81ff0bd4",
  1305 => x"0cd00870",
  1306 => x"8f2a7081",
  1307 => x"06515153",
  1308 => x"72f33872",
  1309 => x"d00c7280",
  1310 => x"c1fc0c02",
  1311 => x"98050d04",
  1312 => x"02e8050d",
  1313 => x"78558056",
  1314 => x"81ff0bd4",
  1315 => x"0cd00870",
  1316 => x"8f2a7081",
  1317 => x"06515153",
  1318 => x"72f33882",
  1319 => x"810bd00c",
  1320 => x"81ff0bd4",
  1321 => x"0c775287",
  1322 => x"fc80d151",
  1323 => x"a2c22d80",
  1324 => x"dbc6df54",
  1325 => x"80c1fc08",
  1326 => x"802e8a38",
  1327 => x"bdfc5186",
  1328 => x"922daa99",
  1329 => x"0481ff0b",
  1330 => x"d40cd408",
  1331 => x"7081ff06",
  1332 => x"51537281",
  1333 => x"fe2e0981",
  1334 => x"069e3880",
  1335 => x"ff53a1f3",
  1336 => x"2d80c1fc",
  1337 => x"08757084",
  1338 => x"05570cff",
  1339 => x"13537280",
  1340 => x"25ec3881",
  1341 => x"56a9fe04",
  1342 => x"ff145473",
  1343 => x"c83881ff",
  1344 => x"0bd40c81",
  1345 => x"ff0bd40c",
  1346 => x"d008708f",
  1347 => x"2a708106",
  1348 => x"51515372",
  1349 => x"f33872d0",
  1350 => x"0c7580c1",
  1351 => x"fc0c0298",
  1352 => x"050d0402",
  1353 => x"f4050d74",
  1354 => x"70882a83",
  1355 => x"fe800670",
  1356 => x"72982a07",
  1357 => x"72882b87",
  1358 => x"fc808006",
  1359 => x"73982b81",
  1360 => x"f00a0671",
  1361 => x"73070780",
  1362 => x"c1fc0c56",
  1363 => x"51535102",
  1364 => x"8c050d04",
  1365 => x"02f8050d",
  1366 => x"028e0580",
  1367 => x"f52d7488",
  1368 => x"2b077083",
  1369 => x"ffff0680",
  1370 => x"c1fc0c51",
  1371 => x"0288050d",
  1372 => x"0402fc05",
  1373 => x"0d725180",
  1374 => x"710c800b",
  1375 => x"84120c02",
  1376 => x"84050d04",
  1377 => x"02f0050d",
  1378 => x"75700884",
  1379 => x"12085353",
  1380 => x"53ff5471",
  1381 => x"712ea838",
  1382 => x"aedb2d84",
  1383 => x"13087084",
  1384 => x"29148811",
  1385 => x"70087081",
  1386 => x"ff068418",
  1387 => x"08811187",
  1388 => x"06841a0c",
  1389 => x"53515551",
  1390 => x"5151aed5",
  1391 => x"2d715473",
  1392 => x"80c1fc0c",
  1393 => x"0290050d",
  1394 => x"0402f805",
  1395 => x"0daedb2d",
  1396 => x"e008708b",
  1397 => x"2a708106",
  1398 => x"51525270",
  1399 => x"802ea138",
  1400 => x"80cbf008",
  1401 => x"70842980",
  1402 => x"cbf80573",
  1403 => x"81ff0671",
  1404 => x"0c515180",
  1405 => x"cbf00881",
  1406 => x"11870680",
  1407 => x"cbf00c51",
  1408 => x"800b80cc",
  1409 => x"980caecd",
  1410 => x"2daed52d",
  1411 => x"0288050d",
  1412 => x"0402fc05",
  1413 => x"0daedb2d",
  1414 => x"810b80cc",
  1415 => x"980caed5",
  1416 => x"2d80cc98",
  1417 => x"085170f9",
  1418 => x"38028405",
  1419 => x"0d0402fc",
  1420 => x"050d80cb",
  1421 => x"f051aaf1",
  1422 => x"2dabc951",
  1423 => x"aec92dad",
  1424 => x"f02d0284",
  1425 => x"050d0402",
  1426 => x"f4050dad",
  1427 => x"d50480c1",
  1428 => x"fc0881f0",
  1429 => x"2e098106",
  1430 => x"8a38810b",
  1431 => x"80c1f00c",
  1432 => x"add50480",
  1433 => x"c1fc0881",
  1434 => x"e02e0981",
  1435 => x"068a3881",
  1436 => x"0b80c1f4",
  1437 => x"0cadd504",
  1438 => x"80c1fc08",
  1439 => x"5280c1f4",
  1440 => x"08802e89",
  1441 => x"3880c1fc",
  1442 => x"08818005",
  1443 => x"5271842c",
  1444 => x"728f0653",
  1445 => x"5380c1f0",
  1446 => x"08802e9a",
  1447 => x"38728429",
  1448 => x"80c1b005",
  1449 => x"72138171",
  1450 => x"2b700973",
  1451 => x"0806730c",
  1452 => x"515353ad",
  1453 => x"c9047284",
  1454 => x"2980c1b0",
  1455 => x"05721383",
  1456 => x"712b7208",
  1457 => x"07720c53",
  1458 => x"53800b80",
  1459 => x"c1f40c80",
  1460 => x"0b80c1f0",
  1461 => x"0c80cbf0",
  1462 => x"51ab842d",
  1463 => x"80c1fc08",
  1464 => x"ff24feea",
  1465 => x"38800b80",
  1466 => x"c1fc0c02",
  1467 => x"8c050d04",
  1468 => x"02f8050d",
  1469 => x"80c1b052",
  1470 => x"8f518072",
  1471 => x"70840554",
  1472 => x"0cff1151",
  1473 => x"708025f2",
  1474 => x"38028805",
  1475 => x"0d0402f0",
  1476 => x"050d7551",
  1477 => x"aedb2d70",
  1478 => x"822cfc06",
  1479 => x"80c1b011",
  1480 => x"72109e06",
  1481 => x"71087072",
  1482 => x"2a708306",
  1483 => x"82742b70",
  1484 => x"09740676",
  1485 => x"0c545156",
  1486 => x"57535153",
  1487 => x"aed52d71",
  1488 => x"80c1fc0c",
  1489 => x"0290050d",
  1490 => x"0471980c",
  1491 => x"04ffb008",
  1492 => x"80c1fc0c",
  1493 => x"04810bff",
  1494 => x"b00c0480",
  1495 => x"0bffb00c",
  1496 => x"0402fc05",
  1497 => x"0d810b80",
  1498 => x"c1f80c81",
  1499 => x"5185812d",
  1500 => x"0284050d",
  1501 => x"0402fc05",
  1502 => x"0d800b80",
  1503 => x"c1f80c80",
  1504 => x"5185812d",
  1505 => x"0284050d",
  1506 => x"0402ec05",
  1507 => x"0d765480",
  1508 => x"52870b88",
  1509 => x"1580f52d",
  1510 => x"56537472",
  1511 => x"248338a0",
  1512 => x"53725182",
  1513 => x"f82d8112",
  1514 => x"8b1580f5",
  1515 => x"2d545272",
  1516 => x"7225de38",
  1517 => x"0294050d",
  1518 => x"0402f005",
  1519 => x"0d80cca8",
  1520 => x"085481f9",
  1521 => x"2d800b80",
  1522 => x"ccac0c73",
  1523 => x"08802e81",
  1524 => x"8638820b",
  1525 => x"80c2900c",
  1526 => x"80ccac08",
  1527 => x"8f0680c2",
  1528 => x"8c0c7308",
  1529 => x"5271832e",
  1530 => x"96387183",
  1531 => x"26893871",
  1532 => x"812eaf38",
  1533 => x"b0c00471",
  1534 => x"852e9f38",
  1535 => x"b0c00488",
  1536 => x"1480f52d",
  1537 => x"841508be",
  1538 => x"8c535452",
  1539 => x"86922d71",
  1540 => x"84291370",
  1541 => x"085252b0",
  1542 => x"c4047351",
  1543 => x"af892db0",
  1544 => x"c00480cc",
  1545 => x"9c088815",
  1546 => x"082c7081",
  1547 => x"06515271",
  1548 => x"802e8738",
  1549 => x"be9051b0",
  1550 => x"bd04be94",
  1551 => x"5186922d",
  1552 => x"84140851",
  1553 => x"86922d80",
  1554 => x"ccac0881",
  1555 => x"0580ccac",
  1556 => x"0c8c1454",
  1557 => x"afcb0402",
  1558 => x"90050d04",
  1559 => x"7180cca8",
  1560 => x"0cafb92d",
  1561 => x"80ccac08",
  1562 => x"ff0580cc",
  1563 => x"b00c0402",
  1564 => x"e8050d80",
  1565 => x"cca80880",
  1566 => x"ccb40857",
  1567 => x"5580f851",
  1568 => x"ae8e2d80",
  1569 => x"c1fc0881",
  1570 => x"2a708106",
  1571 => x"5152719c",
  1572 => x"388751ae",
  1573 => x"8e2d80c1",
  1574 => x"fc08812a",
  1575 => x"70810651",
  1576 => x"5271802e",
  1577 => x"b538b1ac",
  1578 => x"04acc72d",
  1579 => x"8751ae8e",
  1580 => x"2d80c1fc",
  1581 => x"08f338b1",
  1582 => x"bd04acc7",
  1583 => x"2d80f851",
  1584 => x"ae8e2d80",
  1585 => x"c1fc08f2",
  1586 => x"3880c1f8",
  1587 => x"08813270",
  1588 => x"80c1f80c",
  1589 => x"70525285",
  1590 => x"812d800b",
  1591 => x"80cca00c",
  1592 => x"800b80cc",
  1593 => x"a40c80c1",
  1594 => x"f808838d",
  1595 => x"3880da51",
  1596 => x"ae8e2d80",
  1597 => x"c1fc0880",
  1598 => x"2e8c3880",
  1599 => x"cca00881",
  1600 => x"800780cc",
  1601 => x"a00c80d9",
  1602 => x"51ae8e2d",
  1603 => x"80c1fc08",
  1604 => x"802e8c38",
  1605 => x"80cca008",
  1606 => x"80c00780",
  1607 => x"cca00c81",
  1608 => x"9451ae8e",
  1609 => x"2d80c1fc",
  1610 => x"08802e8b",
  1611 => x"3880cca0",
  1612 => x"08900780",
  1613 => x"cca00c81",
  1614 => x"9151ae8e",
  1615 => x"2d80c1fc",
  1616 => x"08802e8b",
  1617 => x"3880cca0",
  1618 => x"08a00780",
  1619 => x"cca00c81",
  1620 => x"f551ae8e",
  1621 => x"2d80c1fc",
  1622 => x"08802e8b",
  1623 => x"3880cca0",
  1624 => x"08810780",
  1625 => x"cca00c81",
  1626 => x"f251ae8e",
  1627 => x"2d80c1fc",
  1628 => x"08802e8b",
  1629 => x"3880cca0",
  1630 => x"08820780",
  1631 => x"cca00c81",
  1632 => x"eb51ae8e",
  1633 => x"2d80c1fc",
  1634 => x"08802e8b",
  1635 => x"3880cca0",
  1636 => x"08840780",
  1637 => x"cca00c81",
  1638 => x"f451ae8e",
  1639 => x"2d80c1fc",
  1640 => x"08802e8b",
  1641 => x"3880cca0",
  1642 => x"08880780",
  1643 => x"cca00c80",
  1644 => x"d851ae8e",
  1645 => x"2d80c1fc",
  1646 => x"08802e8c",
  1647 => x"3880cca4",
  1648 => x"08818007",
  1649 => x"80cca40c",
  1650 => x"9251ae8e",
  1651 => x"2d80c1fc",
  1652 => x"08802e8c",
  1653 => x"3880cca4",
  1654 => x"0880c007",
  1655 => x"80cca40c",
  1656 => x"9451ae8e",
  1657 => x"2d80c1fc",
  1658 => x"08802e8b",
  1659 => x"3880cca4",
  1660 => x"08900780",
  1661 => x"cca40c91",
  1662 => x"51ae8e2d",
  1663 => x"80c1fc08",
  1664 => x"802e8b38",
  1665 => x"80cca408",
  1666 => x"a00780cc",
  1667 => x"a40c9d51",
  1668 => x"ae8e2d80",
  1669 => x"c1fc0880",
  1670 => x"2e8b3880",
  1671 => x"cca40881",
  1672 => x"0780cca4",
  1673 => x"0c9b51ae",
  1674 => x"8e2d80c1",
  1675 => x"fc08802e",
  1676 => x"8b3880cc",
  1677 => x"a4088207",
  1678 => x"80cca40c",
  1679 => x"9c51ae8e",
  1680 => x"2d80c1fc",
  1681 => x"08802e8b",
  1682 => x"3880cca4",
  1683 => x"08840780",
  1684 => x"cca40ca3",
  1685 => x"51ae8e2d",
  1686 => x"80c1fc08",
  1687 => x"802e8b38",
  1688 => x"80cca408",
  1689 => x"880780cc",
  1690 => x"a40c81fd",
  1691 => x"51ae8e2d",
  1692 => x"81fa51ae",
  1693 => x"8e2dbace",
  1694 => x"0481f551",
  1695 => x"ae8e2d80",
  1696 => x"c1fc0881",
  1697 => x"2a708106",
  1698 => x"51527180",
  1699 => x"2eb33880",
  1700 => x"ccb00852",
  1701 => x"71802e8a",
  1702 => x"38ff1280",
  1703 => x"ccb00cb5",
  1704 => x"c10480cc",
  1705 => x"ac081080",
  1706 => x"ccac0805",
  1707 => x"70842916",
  1708 => x"51528812",
  1709 => x"08802e89",
  1710 => x"38ff5188",
  1711 => x"12085271",
  1712 => x"2d81f251",
  1713 => x"ae8e2d80",
  1714 => x"c1fc0881",
  1715 => x"2a708106",
  1716 => x"51527180",
  1717 => x"2eb43880",
  1718 => x"ccac08ff",
  1719 => x"1180ccb0",
  1720 => x"08565353",
  1721 => x"7372258a",
  1722 => x"38811480",
  1723 => x"ccb00cb6",
  1724 => x"8a047210",
  1725 => x"13708429",
  1726 => x"16515288",
  1727 => x"1208802e",
  1728 => x"8938fe51",
  1729 => x"88120852",
  1730 => x"712d81fd",
  1731 => x"51ae8e2d",
  1732 => x"80c1fc08",
  1733 => x"812a7081",
  1734 => x"06515271",
  1735 => x"802eb138",
  1736 => x"80ccb008",
  1737 => x"802e8a38",
  1738 => x"800b80cc",
  1739 => x"b00cb6d0",
  1740 => x"0480ccac",
  1741 => x"081080cc",
  1742 => x"ac080570",
  1743 => x"84291651",
  1744 => x"52881208",
  1745 => x"802e8938",
  1746 => x"fd518812",
  1747 => x"0852712d",
  1748 => x"81fa51ae",
  1749 => x"8e2d80c1",
  1750 => x"fc08812a",
  1751 => x"70810651",
  1752 => x"5271802e",
  1753 => x"b13880cc",
  1754 => x"ac08ff11",
  1755 => x"545280cc",
  1756 => x"b0087325",
  1757 => x"89387280",
  1758 => x"ccb00cb7",
  1759 => x"96047110",
  1760 => x"12708429",
  1761 => x"16515288",
  1762 => x"1208802e",
  1763 => x"8938fc51",
  1764 => x"88120852",
  1765 => x"712d80cc",
  1766 => x"b0087053",
  1767 => x"5473802e",
  1768 => x"8a388c15",
  1769 => x"ff155555",
  1770 => x"b79d0482",
  1771 => x"0b80c290",
  1772 => x"0c718f06",
  1773 => x"80c28c0c",
  1774 => x"81eb51ae",
  1775 => x"8e2d80c1",
  1776 => x"fc08812a",
  1777 => x"70810651",
  1778 => x"5271802e",
  1779 => x"ad387408",
  1780 => x"852e0981",
  1781 => x"06a43888",
  1782 => x"1580f52d",
  1783 => x"ff055271",
  1784 => x"881681b7",
  1785 => x"2d71982b",
  1786 => x"52718025",
  1787 => x"8838800b",
  1788 => x"881681b7",
  1789 => x"2d7451af",
  1790 => x"892d81f4",
  1791 => x"51ae8e2d",
  1792 => x"80c1fc08",
  1793 => x"812a7081",
  1794 => x"06515271",
  1795 => x"802eb338",
  1796 => x"7408852e",
  1797 => x"098106aa",
  1798 => x"38881580",
  1799 => x"f52d8105",
  1800 => x"52718816",
  1801 => x"81b72d71",
  1802 => x"81ff068b",
  1803 => x"1680f52d",
  1804 => x"54527272",
  1805 => x"27873872",
  1806 => x"881681b7",
  1807 => x"2d7451af",
  1808 => x"892d80da",
  1809 => x"51ae8e2d",
  1810 => x"80c1fc08",
  1811 => x"812a7081",
  1812 => x"06515271",
  1813 => x"802e81ad",
  1814 => x"3880cca8",
  1815 => x"0880ccb0",
  1816 => x"08555373",
  1817 => x"802e8a38",
  1818 => x"8c13ff15",
  1819 => x"5553b8e3",
  1820 => x"04720852",
  1821 => x"71822ea6",
  1822 => x"38718226",
  1823 => x"89387181",
  1824 => x"2eaa38ba",
  1825 => x"85047183",
  1826 => x"2eb43871",
  1827 => x"842e0981",
  1828 => x"0680f238",
  1829 => x"88130851",
  1830 => x"b0dc2dba",
  1831 => x"850480cc",
  1832 => x"b0085188",
  1833 => x"13085271",
  1834 => x"2dba8504",
  1835 => x"810b8814",
  1836 => x"082b80cc",
  1837 => x"9c083280",
  1838 => x"cc9c0cb9",
  1839 => x"d9048813",
  1840 => x"80f52d81",
  1841 => x"058b1480",
  1842 => x"f52d5354",
  1843 => x"71742483",
  1844 => x"38805473",
  1845 => x"881481b7",
  1846 => x"2dafb92d",
  1847 => x"ba850475",
  1848 => x"08802ea4",
  1849 => x"38750851",
  1850 => x"ae8e2d80",
  1851 => x"c1fc0881",
  1852 => x"06527180",
  1853 => x"2e8c3880",
  1854 => x"ccb00851",
  1855 => x"84160852",
  1856 => x"712d8816",
  1857 => x"5675d838",
  1858 => x"8054800b",
  1859 => x"80c2900c",
  1860 => x"738f0680",
  1861 => x"c28c0ca0",
  1862 => x"527380cc",
  1863 => x"b0082e09",
  1864 => x"81069938",
  1865 => x"80ccac08",
  1866 => x"ff057432",
  1867 => x"70098105",
  1868 => x"7072079f",
  1869 => x"2a917131",
  1870 => x"51515353",
  1871 => x"715182f8",
  1872 => x"2d811454",
  1873 => x"8e7425c2",
  1874 => x"3880c1f8",
  1875 => x"08527180",
  1876 => x"c1fc0c02",
  1877 => x"98050d04",
  1878 => x"00ffffff",
  1879 => x"ff00ffff",
  1880 => x"ffff00ff",
  1881 => x"ffffff00",
  1882 => x"4f4b0000",
  1883 => x"52657365",
  1884 => x"74000000",
  1885 => x"53617665",
  1886 => x"20736574",
  1887 => x"74696e67",
  1888 => x"73000000",
  1889 => x"5363616e",
  1890 => x"6c696e65",
  1891 => x"73000000",
  1892 => x"41756469",
  1893 => x"6f20566f",
  1894 => x"6c756d65",
  1895 => x"00000000",
  1896 => x"4c6f6164",
  1897 => x"20524f4d",
  1898 => x"20100000",
  1899 => x"45786974",
  1900 => x"00000000",
  1901 => x"464d2064",
  1902 => x"69736162",
  1903 => x"6c650000",
  1904 => x"464d2065",
  1905 => x"6e61626c",
  1906 => x"65000000",
  1907 => x"50534720",
  1908 => x"64697361",
  1909 => x"626c6500",
  1910 => x"50534720",
  1911 => x"656e6162",
  1912 => x"6c650000",
  1913 => x"4a6f7973",
  1914 => x"7469636b",
  1915 => x"20737761",
  1916 => x"70000000",
  1917 => x"4a6f7973",
  1918 => x"7469636b",
  1919 => x"206e6f72",
  1920 => x"6d616c00",
  1921 => x"56474120",
  1922 => x"2d203331",
  1923 => x"4b487a00",
  1924 => x"5456202d",
  1925 => x"2031354b",
  1926 => x"487a0000",
  1927 => x"4261636b",
  1928 => x"00000000",
  1929 => x"4c6f6164",
  1930 => x"20457272",
  1931 => x"6f722100",
  1932 => x"46504741",
  1933 => x"47454e20",
  1934 => x"43464700",
  1935 => x"496e6974",
  1936 => x"69616c69",
  1937 => x"7a696e67",
  1938 => x"20534420",
  1939 => x"63617264",
  1940 => x"0a000000",
  1941 => x"424f4f54",
  1942 => x"20202020",
  1943 => x"47454e00",
  1944 => x"43617264",
  1945 => x"20696e69",
  1946 => x"74206661",
  1947 => x"696c6564",
  1948 => x"0a000000",
  1949 => x"4d425220",
  1950 => x"6661696c",
  1951 => x"0a000000",
  1952 => x"46415431",
  1953 => x"36202020",
  1954 => x"00000000",
  1955 => x"46415433",
  1956 => x"32202020",
  1957 => x"00000000",
  1958 => x"4e6f2070",
  1959 => x"61727469",
  1960 => x"74696f6e",
  1961 => x"20736967",
  1962 => x"0a000000",
  1963 => x"42616420",
  1964 => x"70617274",
  1965 => x"0a000000",
  1966 => x"53444843",
  1967 => x"20657272",
  1968 => x"6f72210a",
  1969 => x"00000000",
  1970 => x"53442069",
  1971 => x"6e69742e",
  1972 => x"2e2e0a00",
  1973 => x"53442063",
  1974 => x"61726420",
  1975 => x"72657365",
  1976 => x"74206661",
  1977 => x"696c6564",
  1978 => x"210a0000",
  1979 => x"57726974",
  1980 => x"65206661",
  1981 => x"696c6564",
  1982 => x"0a000000",
  1983 => x"52656164",
  1984 => x"20666169",
  1985 => x"6c65640a",
  1986 => x"00000000",
  1987 => x"16200000",
  1988 => x"14200000",
  1989 => x"15200000",
  1990 => x"00000002",
  1991 => x"00000000",
  1992 => x"00000002",
  1993 => x"00001d6c",
  1994 => x"000004ff",
  1995 => x"00000002",
  1996 => x"00001d74",
  1997 => x"000003c4",
  1998 => x"00000003",
  1999 => x"00001fbc",
  2000 => x"00000002",
  2001 => x"00000001",
  2002 => x"00001d84",
  2003 => x"00000001",
  2004 => x"00000003",
  2005 => x"00001fb4",
  2006 => x"00000002",
  2007 => x"00000005",
  2008 => x"00001d90",
  2009 => x"00000007",
  2010 => x"00000003",
  2011 => x"00001fac",
  2012 => x"00000002",
  2013 => x"00000003",
  2014 => x"00001fa4",
  2015 => x"00000002",
  2016 => x"00000002",
  2017 => x"00001da0",
  2018 => x"000007d3",
  2019 => x"00000002",
  2020 => x"00001dac",
  2021 => x"00001775",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00001db4",
  2026 => x"00001dc0",
  2027 => x"00001dcc",
  2028 => x"00001dd8",
  2029 => x"00001de4",
  2030 => x"00001df4",
  2031 => x"00001e04",
  2032 => x"00001e10",
  2033 => x"00000002",
  2034 => x"00002128",
  2035 => x"00000591",
  2036 => x"00000002",
  2037 => x"00002146",
  2038 => x"00000591",
  2039 => x"00000002",
  2040 => x"00002164",
  2041 => x"00000591",
  2042 => x"00000002",
  2043 => x"00002182",
  2044 => x"00000591",
  2045 => x"00000002",
  2046 => x"000021a0",
  2047 => x"00000591",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

