-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b0bbe",
     9 => x"88080b0b",
    10 => x"0bbe8c08",
    11 => x"0b0b0bbe",
    12 => x"90080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"be900c0b",
    16 => x"0b0bbe8c",
    17 => x"0c0b0b0b",
    18 => x"be880c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb7f4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"be887080",
    57 => x"c8c8278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"518fe204",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbe980c",
    65 => x"9f0bbe9c",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"be9c08ff",
    69 => x"05be9c0c",
    70 => x"be9c0880",
    71 => x"25eb38be",
    72 => x"9808ff05",
    73 => x"be980cbe",
    74 => x"98088025",
    75 => x"d7380284",
    76 => x"050d0402",
    77 => x"f0050df8",
    78 => x"8053f8a0",
    79 => x"5483bf52",
    80 => x"73708105",
    81 => x"55335170",
    82 => x"73708105",
    83 => x"5534ff12",
    84 => x"52718025",
    85 => x"eb38fbc0",
    86 => x"539f52a0",
    87 => x"73708105",
    88 => x"5534ff12",
    89 => x"52718025",
    90 => x"f2380290",
    91 => x"050d0402",
    92 => x"f4050d74",
    93 => x"538e0bbe",
    94 => x"9808258f",
    95 => x"3882b32d",
    96 => x"be9808ff",
    97 => x"05be980c",
    98 => x"82f504be",
    99 => x"9808be9c",
   100 => x"08535172",
   101 => x"8a2e0981",
   102 => x"06b73871",
   103 => x"51719f24",
   104 => x"a038be98",
   105 => x"08a02911",
   106 => x"f8801151",
   107 => x"51a07134",
   108 => x"be9c0881",
   109 => x"05be9c0c",
   110 => x"be9c0851",
   111 => x"9f7125e2",
   112 => x"38800bbe",
   113 => x"9c0cbe98",
   114 => x"088105be",
   115 => x"980c83e5",
   116 => x"0470a029",
   117 => x"12f88011",
   118 => x"51517271",
   119 => x"34be9c08",
   120 => x"8105be9c",
   121 => x"0cbe9c08",
   122 => x"a02e0981",
   123 => x"068e3880",
   124 => x"0bbe9c0c",
   125 => x"be980881",
   126 => x"05be980c",
   127 => x"028c050d",
   128 => x"0402e805",
   129 => x"0d777956",
   130 => x"56880bfc",
   131 => x"1677712c",
   132 => x"8f065452",
   133 => x"54805372",
   134 => x"72259538",
   135 => x"7153fbe0",
   136 => x"14518771",
   137 => x"348114ff",
   138 => x"14545472",
   139 => x"f1387153",
   140 => x"f9157671",
   141 => x"2c870653",
   142 => x"5171802e",
   143 => x"8b38fbe0",
   144 => x"14517171",
   145 => x"34811454",
   146 => x"728e2495",
   147 => x"388f7331",
   148 => x"53fbe014",
   149 => x"51a07134",
   150 => x"8114ff14",
   151 => x"545472f1",
   152 => x"38029805",
   153 => x"0d0402ec",
   154 => x"050d800b",
   155 => x"bea00cf6",
   156 => x"8c08f690",
   157 => x"0871882c",
   158 => x"565481ff",
   159 => x"06527372",
   160 => x"25883871",
   161 => x"54820bbe",
   162 => x"a00c7288",
   163 => x"2c7381ff",
   164 => x"06545574",
   165 => x"73258b38",
   166 => x"72bea008",
   167 => x"8407bea0",
   168 => x"0c557384",
   169 => x"2b87e871",
   170 => x"25837131",
   171 => x"700b0b0b",
   172 => x"baf40c81",
   173 => x"712bf688",
   174 => x"0cfea413",
   175 => x"ff122c78",
   176 => x"8829ff94",
   177 => x"0570812c",
   178 => x"bea00852",
   179 => x"58525551",
   180 => x"52547680",
   181 => x"2e853870",
   182 => x"81075170",
   183 => x"f6940c71",
   184 => x"098105f6",
   185 => x"800c7209",
   186 => x"8105f684",
   187 => x"0c029405",
   188 => x"0d0402f4",
   189 => x"050d7453",
   190 => x"72708105",
   191 => x"5480f52d",
   192 => x"5271802e",
   193 => x"89387151",
   194 => x"82ef2d85",
   195 => x"f804028c",
   196 => x"050d0402",
   197 => x"f4050d74",
   198 => x"70820680",
   199 => x"c8ac0cbb",
   200 => x"90718106",
   201 => x"54545171",
   202 => x"881481b7",
   203 => x"2d70822a",
   204 => x"70810651",
   205 => x"5170a014",
   206 => x"81b72d70",
   207 => x"be880c02",
   208 => x"8c050d04",
   209 => x"02f8050d",
   210 => x"b98c52be",
   211 => x"a4519ccc",
   212 => x"2dbe8808",
   213 => x"802ea138",
   214 => x"80c1c052",
   215 => x"bea4519f",
   216 => x"8d2d80c1",
   217 => x"c008beb0",
   218 => x"0c80c1c0",
   219 => x"08fec00c",
   220 => x"80c1c008",
   221 => x"5186932d",
   222 => x"0288050d",
   223 => x"0402f005",
   224 => x"0d805192",
   225 => x"9b2db98c",
   226 => x"52bea451",
   227 => x"9ccc2dbe",
   228 => x"8808802e",
   229 => x"a838beb0",
   230 => x"0880c1c0",
   231 => x"0c80c1c4",
   232 => x"5480fd53",
   233 => x"80747084",
   234 => x"05560cff",
   235 => x"13537280",
   236 => x"25f23880",
   237 => x"c1c052be",
   238 => x"a4519fb6",
   239 => x"2d029005",
   240 => x"0d0402d4",
   241 => x"050dbeb0",
   242 => x"08fec00c",
   243 => x"810bfec4",
   244 => x"0c840bfe",
   245 => x"c40c7c52",
   246 => x"bea4519c",
   247 => x"cc2dbe88",
   248 => x"0853be88",
   249 => x"08802e81",
   250 => x"ce38bea8",
   251 => x"0856800b",
   252 => x"ff175859",
   253 => x"76792e8b",
   254 => x"38811977",
   255 => x"812a5859",
   256 => x"76f738f7",
   257 => x"19769fff",
   258 => x"06545972",
   259 => x"802e8b38",
   260 => x"fc8016be",
   261 => x"a452569e",
   262 => x"df2d75b0",
   263 => x"80802e09",
   264 => x"81068938",
   265 => x"820bfedc",
   266 => x"0c88c304",
   267 => x"75988080",
   268 => x"2e098106",
   269 => x"8938810b",
   270 => x"fedc0c88",
   271 => x"c304800b",
   272 => x"fedc0c81",
   273 => x"5b807625",
   274 => x"80eb3878",
   275 => x"52765184",
   276 => x"812d80c1",
   277 => x"c052bea4",
   278 => x"519f8d2d",
   279 => x"be880880",
   280 => x"2ebc3880",
   281 => x"c1c05a83",
   282 => x"fc587970",
   283 => x"84055b08",
   284 => x"7083fe80",
   285 => x"0671882b",
   286 => x"83fe8006",
   287 => x"71882a07",
   288 => x"72882a83",
   289 => x"fe800673",
   290 => x"982a07fe",
   291 => x"c80cfec8",
   292 => x"0c56fc19",
   293 => x"59537780",
   294 => x"25d03889",
   295 => x"a504be88",
   296 => x"085b8480",
   297 => x"56bea451",
   298 => x"9edf2dfc",
   299 => x"80168118",
   300 => x"585688c5",
   301 => x"047a5372",
   302 => x"be880c02",
   303 => x"ac050d04",
   304 => x"02fc050d",
   305 => x"acb32dfe",
   306 => x"c4518171",
   307 => x"0c82710c",
   308 => x"0284050d",
   309 => x"0402f405",
   310 => x"0d747678",
   311 => x"53545280",
   312 => x"71259738",
   313 => x"72708105",
   314 => x"5480f52d",
   315 => x"72708105",
   316 => x"5481b72d",
   317 => x"ff115170",
   318 => x"eb388072",
   319 => x"81b72d02",
   320 => x"8c050d04",
   321 => x"02e8050d",
   322 => x"77568070",
   323 => x"56547376",
   324 => x"24b33880",
   325 => x"c7d00874",
   326 => x"2eab3873",
   327 => x"519a952d",
   328 => x"be8808be",
   329 => x"88080981",
   330 => x"0570be88",
   331 => x"08079f2a",
   332 => x"77058117",
   333 => x"57575353",
   334 => x"74762489",
   335 => x"3880c7d0",
   336 => x"087426d7",
   337 => x"3872be88",
   338 => x"0c029805",
   339 => x"0d0402f4",
   340 => x"050dbdb4",
   341 => x"0815518a",
   342 => x"842dbe88",
   343 => x"08802e95",
   344 => x"388b53be",
   345 => x"88085280",
   346 => x"c5c05189",
   347 => x"d52d80c5",
   348 => x"c05187c2",
   349 => x"2dbaf851",
   350 => x"ae972dac",
   351 => x"b32d8051",
   352 => x"84e62d02",
   353 => x"8c050d04",
   354 => x"02dc050d",
   355 => x"80705a55",
   356 => x"74bdb408",
   357 => x"25b13880",
   358 => x"c7d00875",
   359 => x"2ea93878",
   360 => x"519a952d",
   361 => x"be880809",
   362 => x"810570be",
   363 => x"8808079f",
   364 => x"2a760581",
   365 => x"1b5b5654",
   366 => x"74bdb408",
   367 => x"25893880",
   368 => x"c7d00879",
   369 => x"26d93880",
   370 => x"557880c7",
   371 => x"d0082781",
   372 => x"d0387851",
   373 => x"9a952dbe",
   374 => x"8808802e",
   375 => x"81a538be",
   376 => x"88088b05",
   377 => x"80f52d70",
   378 => x"842a7081",
   379 => x"06771078",
   380 => x"842b80c5",
   381 => x"c00b80f5",
   382 => x"2d5c5c53",
   383 => x"51555673",
   384 => x"802e80c7",
   385 => x"38741682",
   386 => x"2b8dc40b",
   387 => x"bc88120c",
   388 => x"54777531",
   389 => x"10beb811",
   390 => x"55569074",
   391 => x"70810556",
   392 => x"81b72da0",
   393 => x"7481b72d",
   394 => x"7681ff06",
   395 => x"81165854",
   396 => x"73802e8a",
   397 => x"389c5380",
   398 => x"c5c0528c",
   399 => x"c4048b53",
   400 => x"be880852",
   401 => x"beba1651",
   402 => x"8cfb0474",
   403 => x"16822b8a",
   404 => x"ce0bbc88",
   405 => x"120c5476",
   406 => x"81ff0681",
   407 => x"16585473",
   408 => x"802e8a38",
   409 => x"9c5380c5",
   410 => x"c0528cf3",
   411 => x"048b53be",
   412 => x"88085277",
   413 => x"753110be",
   414 => x"b8055176",
   415 => x"5589d52d",
   416 => x"8d960474",
   417 => x"90297531",
   418 => x"7010beb8",
   419 => x"055154be",
   420 => x"88087481",
   421 => x"b72d8119",
   422 => x"59748b24",
   423 => x"a2388bc9",
   424 => x"04749029",
   425 => x"75317010",
   426 => x"beb8058c",
   427 => x"77315751",
   428 => x"54807481",
   429 => x"b72d9e14",
   430 => x"ff165654",
   431 => x"74f33802",
   432 => x"a4050d04",
   433 => x"02fc050d",
   434 => x"bdb40813",
   435 => x"518a842d",
   436 => x"be880880",
   437 => x"2e8838be",
   438 => x"88085192",
   439 => x"9b2d800b",
   440 => x"bdb40c8b",
   441 => x"882dacf6",
   442 => x"2d028405",
   443 => x"0d0402fc",
   444 => x"050d7251",
   445 => x"70fd2ead",
   446 => x"3870fd24",
   447 => x"8a3870fc",
   448 => x"2e80c438",
   449 => x"8ecf0470",
   450 => x"fe2eb138",
   451 => x"70ff2e09",
   452 => x"8106bc38",
   453 => x"bdb40851",
   454 => x"70802eb3",
   455 => x"38ff11bd",
   456 => x"b40c8ecf",
   457 => x"04bdb408",
   458 => x"f00570bd",
   459 => x"b40c5170",
   460 => x"80259c38",
   461 => x"800bbdb4",
   462 => x"0c8ecf04",
   463 => x"bdb40881",
   464 => x"05bdb40c",
   465 => x"8ecf04bd",
   466 => x"b4089005",
   467 => x"bdb40c8b",
   468 => x"882dacf6",
   469 => x"2d028405",
   470 => x"0d0402fc",
   471 => x"050dbeb0",
   472 => x"08fb06be",
   473 => x"b00c7251",
   474 => x"8ace2d02",
   475 => x"84050d04",
   476 => x"02fc050d",
   477 => x"beb00884",
   478 => x"07beb00c",
   479 => x"72518ace",
   480 => x"2d028405",
   481 => x"0d0402fc",
   482 => x"050d800b",
   483 => x"bdb40c8b",
   484 => x"882dbc80",
   485 => x"51ae972d",
   486 => x"bbe851ae",
   487 => x"aa2d0284",
   488 => x"050d0402",
   489 => x"f8050d80",
   490 => x"c8ac0882",
   491 => x"06bb980b",
   492 => x"80f52d52",
   493 => x"5270802e",
   494 => x"85387181",
   495 => x"0752bbb0",
   496 => x"0b80f52d",
   497 => x"5170802e",
   498 => x"85387184",
   499 => x"0752beb4",
   500 => x"08802e85",
   501 => x"38719007",
   502 => x"5271be88",
   503 => x"0c028805",
   504 => x"0d0402f4",
   505 => x"050d810b",
   506 => x"beb40c90",
   507 => x"5186932d",
   508 => x"810bfec4",
   509 => x"0c900bfe",
   510 => x"c00c840b",
   511 => x"fec40c83",
   512 => x"0bfecc0c",
   513 => x"a9ff2dac",
   514 => x"942da9e2",
   515 => x"2da9e22d",
   516 => x"81f82d81",
   517 => x"5184e62d",
   518 => x"a9e22da9",
   519 => x"e22d8151",
   520 => x"84e62db9",
   521 => x"985185f2",
   522 => x"2d8452a3",
   523 => x"ed2d93bc",
   524 => x"2dbe8808",
   525 => x"802e8638",
   526 => x"fe5290c5",
   527 => x"04ff1252",
   528 => x"718024e7",
   529 => x"3871802e",
   530 => x"81833886",
   531 => x"c42db9b0",
   532 => x"5187c22d",
   533 => x"be880880",
   534 => x"2e8f38ba",
   535 => x"f851ae97",
   536 => x"2d805184",
   537 => x"e62d90f3",
   538 => x"04be8808",
   539 => x"518f862d",
   540 => x"aca02daa",
   541 => x"982daeb0",
   542 => x"2dbe8808",
   543 => x"80c8b008",
   544 => x"882b80c8",
   545 => x"b40807fe",
   546 => x"d80c538f",
   547 => x"a32dbe88",
   548 => x"08beb008",
   549 => x"2ea238be",
   550 => x"8808beb0",
   551 => x"0cbe8808",
   552 => x"fec00c84",
   553 => x"52725184",
   554 => x"e62da9e2",
   555 => x"2da9e22d",
   556 => x"ff125271",
   557 => x"8025ee38",
   558 => x"72802e89",
   559 => x"388a0bfe",
   560 => x"c40c90f3",
   561 => x"04820bfe",
   562 => x"c40c90f3",
   563 => x"04b9bc51",
   564 => x"85f22d80",
   565 => x"0bbe880c",
   566 => x"028c050d",
   567 => x"0402e805",
   568 => x"0d77797b",
   569 => x"58555580",
   570 => x"53727625",
   571 => x"a3387470",
   572 => x"81055680",
   573 => x"f52d7470",
   574 => x"81055680",
   575 => x"f52d5252",
   576 => x"71712e86",
   577 => x"38815192",
   578 => x"92048113",
   579 => x"5391e904",
   580 => x"805170be",
   581 => x"880c0298",
   582 => x"050d0402",
   583 => x"ec050d76",
   584 => x"5574802e",
   585 => x"be389a15",
   586 => x"80e02d51",
   587 => x"a8a72dbe",
   588 => x"8808be88",
   589 => x"0880c7f0",
   590 => x"0cbe8808",
   591 => x"545480c7",
   592 => x"cc08802e",
   593 => x"99389415",
   594 => x"80e02d51",
   595 => x"a8a72dbe",
   596 => x"8808902b",
   597 => x"83fff00a",
   598 => x"06707507",
   599 => x"51537280",
   600 => x"c7f00c80",
   601 => x"c7f00853",
   602 => x"72802e9d",
   603 => x"3880c7c4",
   604 => x"08fe1471",
   605 => x"2980c7d8",
   606 => x"080580c7",
   607 => x"f40c7084",
   608 => x"2b80c7d0",
   609 => x"0c5493b7",
   610 => x"0480c7dc",
   611 => x"0880c7f0",
   612 => x"0c80c7e0",
   613 => x"0880c7f4",
   614 => x"0c80c7cc",
   615 => x"08802e8b",
   616 => x"3880c7c4",
   617 => x"08842b53",
   618 => x"93b20480",
   619 => x"c7e40884",
   620 => x"2b537280",
   621 => x"c7d00c02",
   622 => x"94050d04",
   623 => x"02d8050d",
   624 => x"800b80c7",
   625 => x"cc0c80c1",
   626 => x"c0528051",
   627 => x"a6d72dbe",
   628 => x"880854be",
   629 => x"88088c38",
   630 => x"b9d05185",
   631 => x"f22d7355",
   632 => x"99980480",
   633 => x"56810b80",
   634 => x"c7f80c88",
   635 => x"53b9dc52",
   636 => x"80c1f651",
   637 => x"91dd2dbe",
   638 => x"8808762e",
   639 => x"09810688",
   640 => x"38be8808",
   641 => x"80c7f80c",
   642 => x"8853b9e8",
   643 => x"5280c292",
   644 => x"5191dd2d",
   645 => x"be880888",
   646 => x"38be8808",
   647 => x"80c7f80c",
   648 => x"80c7f808",
   649 => x"802e80fd",
   650 => x"3880c586",
   651 => x"0b80f52d",
   652 => x"80c5870b",
   653 => x"80f52d71",
   654 => x"982b7190",
   655 => x"2b0780c5",
   656 => x"880b80f5",
   657 => x"2d70882b",
   658 => x"720780c5",
   659 => x"890b80f5",
   660 => x"2d710780",
   661 => x"c5be0b80",
   662 => x"f52d80c5",
   663 => x"bf0b80f5",
   664 => x"2d71882b",
   665 => x"07535f54",
   666 => x"525a5657",
   667 => x"557381ab",
   668 => x"aa2e0981",
   669 => x"068d3875",
   670 => x"51a7f72d",
   671 => x"be880856",
   672 => x"95900473",
   673 => x"82d4d52e",
   674 => x"8738b9f4",
   675 => x"5195d504",
   676 => x"80c1c052",
   677 => x"7551a6d7",
   678 => x"2dbe8808",
   679 => x"55be8808",
   680 => x"802e83f4",
   681 => x"388853b9",
   682 => x"e85280c2",
   683 => x"925191dd",
   684 => x"2dbe8808",
   685 => x"8a38810b",
   686 => x"80c7cc0c",
   687 => x"95db0488",
   688 => x"53b9dc52",
   689 => x"80c1f651",
   690 => x"91dd2dbe",
   691 => x"8808802e",
   692 => x"8a38ba88",
   693 => x"5185f22d",
   694 => x"96ba0480",
   695 => x"c5be0b80",
   696 => x"f52d5473",
   697 => x"80d52e09",
   698 => x"810680ce",
   699 => x"3880c5bf",
   700 => x"0b80f52d",
   701 => x"547381aa",
   702 => x"2e098106",
   703 => x"bd38800b",
   704 => x"80c1c00b",
   705 => x"80f52d56",
   706 => x"547481e9",
   707 => x"2e833881",
   708 => x"547481eb",
   709 => x"2e8c3880",
   710 => x"5573752e",
   711 => x"09810682",
   712 => x"f73880c1",
   713 => x"cb0b80f5",
   714 => x"2d55748e",
   715 => x"3880c1cc",
   716 => x"0b80f52d",
   717 => x"5473822e",
   718 => x"86388055",
   719 => x"99980480",
   720 => x"c1cd0b80",
   721 => x"f52d7080",
   722 => x"c7c40cff",
   723 => x"0580c7c8",
   724 => x"0c80c1ce",
   725 => x"0b80f52d",
   726 => x"80c1cf0b",
   727 => x"80f52d58",
   728 => x"76057782",
   729 => x"80290570",
   730 => x"80c7d40c",
   731 => x"80c1d00b",
   732 => x"80f52d70",
   733 => x"80c7e80c",
   734 => x"80c7cc08",
   735 => x"59575876",
   736 => x"802e81b5",
   737 => x"388853b9",
   738 => x"e85280c2",
   739 => x"925191dd",
   740 => x"2dbe8808",
   741 => x"82823880",
   742 => x"c7c40870",
   743 => x"842b80c7",
   744 => x"d00c7080",
   745 => x"c7e40c80",
   746 => x"c1e50b80",
   747 => x"f52d80c1",
   748 => x"e40b80f5",
   749 => x"2d718280",
   750 => x"290580c1",
   751 => x"e60b80f5",
   752 => x"2d708480",
   753 => x"80291280",
   754 => x"c1e70b80",
   755 => x"f52d7081",
   756 => x"800a2912",
   757 => x"7080c7ec",
   758 => x"0c80c7e8",
   759 => x"08712980",
   760 => x"c7d40805",
   761 => x"7080c7d8",
   762 => x"0c80c1ed",
   763 => x"0b80f52d",
   764 => x"80c1ec0b",
   765 => x"80f52d71",
   766 => x"82802905",
   767 => x"80c1ee0b",
   768 => x"80f52d70",
   769 => x"84808029",
   770 => x"1280c1ef",
   771 => x"0b80f52d",
   772 => x"70982b81",
   773 => x"f00a0672",
   774 => x"057080c7",
   775 => x"dc0cfe11",
   776 => x"7e297705",
   777 => x"80c7e00c",
   778 => x"52595243",
   779 => x"545e5152",
   780 => x"59525d57",
   781 => x"59579991",
   782 => x"0480c1d2",
   783 => x"0b80f52d",
   784 => x"80c1d10b",
   785 => x"80f52d71",
   786 => x"82802905",
   787 => x"7080c7d0",
   788 => x"0c70a029",
   789 => x"83ff0570",
   790 => x"892a7080",
   791 => x"c7e40c80",
   792 => x"c1d70b80",
   793 => x"f52d80c1",
   794 => x"d60b80f5",
   795 => x"2d718280",
   796 => x"29057080",
   797 => x"c7ec0c7b",
   798 => x"71291e70",
   799 => x"80c7e00c",
   800 => x"7d80c7dc",
   801 => x"0c730580",
   802 => x"c7d80c55",
   803 => x"5e515155",
   804 => x"55805192",
   805 => x"9b2d8155",
   806 => x"74be880c",
   807 => x"02a8050d",
   808 => x"0402ec05",
   809 => x"0d767087",
   810 => x"2c7180ff",
   811 => x"06555654",
   812 => x"80c7cc08",
   813 => x"8a387388",
   814 => x"2c7481ff",
   815 => x"06545580",
   816 => x"c1c05280",
   817 => x"c7d40815",
   818 => x"51a6d72d",
   819 => x"be880854",
   820 => x"be880880",
   821 => x"2eb63880",
   822 => x"c7cc0880",
   823 => x"2e993872",
   824 => x"842980c1",
   825 => x"c0057008",
   826 => x"5253a7f7",
   827 => x"2dbe8808",
   828 => x"f00a0653",
   829 => x"9a8a0472",
   830 => x"1080c1c0",
   831 => x"057080e0",
   832 => x"2d5253a8",
   833 => x"a72dbe88",
   834 => x"08537254",
   835 => x"73be880c",
   836 => x"0294050d",
   837 => x"0402e005",
   838 => x"0d797084",
   839 => x"2c80c7f4",
   840 => x"0805718f",
   841 => x"06525553",
   842 => x"728a3880",
   843 => x"c1c05273",
   844 => x"51a6d72d",
   845 => x"72a02980",
   846 => x"c1c00554",
   847 => x"807480f5",
   848 => x"2d565374",
   849 => x"732e8338",
   850 => x"81537481",
   851 => x"e52e81f1",
   852 => x"38817074",
   853 => x"06545872",
   854 => x"802e81e5",
   855 => x"388b1480",
   856 => x"f52d7083",
   857 => x"2a790658",
   858 => x"56769938",
   859 => x"bdb80853",
   860 => x"72893872",
   861 => x"80c5c00b",
   862 => x"81b72d76",
   863 => x"bdb80c73",
   864 => x"539cc304",
   865 => x"758f2e09",
   866 => x"810681b5",
   867 => x"38749f06",
   868 => x"8d2980c5",
   869 => x"b3115153",
   870 => x"811480f5",
   871 => x"2d737081",
   872 => x"055581b7",
   873 => x"2d831480",
   874 => x"f52d7370",
   875 => x"81055581",
   876 => x"b72d8514",
   877 => x"80f52d73",
   878 => x"70810555",
   879 => x"81b72d87",
   880 => x"1480f52d",
   881 => x"73708105",
   882 => x"5581b72d",
   883 => x"891480f5",
   884 => x"2d737081",
   885 => x"055581b7",
   886 => x"2d8e1480",
   887 => x"f52d7370",
   888 => x"81055581",
   889 => x"b72d9014",
   890 => x"80f52d73",
   891 => x"70810555",
   892 => x"81b72d92",
   893 => x"1480f52d",
   894 => x"73708105",
   895 => x"5581b72d",
   896 => x"941480f5",
   897 => x"2d737081",
   898 => x"055581b7",
   899 => x"2d961480",
   900 => x"f52d7370",
   901 => x"81055581",
   902 => x"b72d9814",
   903 => x"80f52d73",
   904 => x"70810555",
   905 => x"81b72d9c",
   906 => x"1480f52d",
   907 => x"73708105",
   908 => x"5581b72d",
   909 => x"9e1480f5",
   910 => x"2d7381b7",
   911 => x"2d77bdb8",
   912 => x"0c805372",
   913 => x"be880c02",
   914 => x"a0050d04",
   915 => x"02cc050d",
   916 => x"7e605e5a",
   917 => x"800b80c7",
   918 => x"f00880c7",
   919 => x"f408595c",
   920 => x"56805880",
   921 => x"c7d00878",
   922 => x"2e81b238",
   923 => x"778f06a0",
   924 => x"17575473",
   925 => x"913880c1",
   926 => x"c0527651",
   927 => x"811757a6",
   928 => x"d72d80c1",
   929 => x"c0568076",
   930 => x"80f52d56",
   931 => x"5474742e",
   932 => x"83388154",
   933 => x"7481e52e",
   934 => x"80f73881",
   935 => x"70750655",
   936 => x"5c73802e",
   937 => x"80eb388b",
   938 => x"1680f52d",
   939 => x"98065978",
   940 => x"80df388b",
   941 => x"537c5275",
   942 => x"5191dd2d",
   943 => x"be880880",
   944 => x"d0389c16",
   945 => x"0851a7f7",
   946 => x"2dbe8808",
   947 => x"841b0c9a",
   948 => x"1680e02d",
   949 => x"51a8a72d",
   950 => x"be8808be",
   951 => x"8808881c",
   952 => x"0cbe8808",
   953 => x"555580c7",
   954 => x"cc08802e",
   955 => x"98389416",
   956 => x"80e02d51",
   957 => x"a8a72dbe",
   958 => x"8808902b",
   959 => x"83fff00a",
   960 => x"06701651",
   961 => x"5473881b",
   962 => x"0c787a0c",
   963 => x"7b549ed6",
   964 => x"04811858",
   965 => x"80c7d008",
   966 => x"7826fed0",
   967 => x"3880c7cc",
   968 => x"08802eb0",
   969 => x"387a5199",
   970 => x"a12dbe88",
   971 => x"08be8808",
   972 => x"80ffffff",
   973 => x"f806555b",
   974 => x"7380ffff",
   975 => x"fff82e94",
   976 => x"38be8808",
   977 => x"fe0580c7",
   978 => x"c4082980",
   979 => x"c7d80805",
   980 => x"579ce104",
   981 => x"805473be",
   982 => x"880c02b4",
   983 => x"050d0402",
   984 => x"f4050d74",
   985 => x"70088105",
   986 => x"710c7008",
   987 => x"80c7c808",
   988 => x"06535371",
   989 => x"8e388813",
   990 => x"085199a1",
   991 => x"2dbe8808",
   992 => x"88140c81",
   993 => x"0bbe880c",
   994 => x"028c050d",
   995 => x"0402f005",
   996 => x"0d758811",
   997 => x"08fe0580",
   998 => x"c7c40829",
   999 => x"80c7d808",
  1000 => x"11720880",
  1001 => x"c7c80806",
  1002 => x"05795553",
  1003 => x"5454a6d7",
  1004 => x"2d029005",
  1005 => x"0d0402f0",
  1006 => x"050d7588",
  1007 => x"1108fe05",
  1008 => x"80c7c408",
  1009 => x"2980c7d8",
  1010 => x"08117208",
  1011 => x"80c7c808",
  1012 => x"06057955",
  1013 => x"535454a5",
  1014 => x"972d0290",
  1015 => x"050d0402",
  1016 => x"f4050dd4",
  1017 => x"5281ff72",
  1018 => x"0c710853",
  1019 => x"81ff720c",
  1020 => x"72882b83",
  1021 => x"fe800672",
  1022 => x"087081ff",
  1023 => x"06515253",
  1024 => x"81ff720c",
  1025 => x"72710788",
  1026 => x"2b720870",
  1027 => x"81ff0651",
  1028 => x"525381ff",
  1029 => x"720c7271",
  1030 => x"07882b72",
  1031 => x"087081ff",
  1032 => x"067207be",
  1033 => x"880c5253",
  1034 => x"028c050d",
  1035 => x"0402f405",
  1036 => x"0d747671",
  1037 => x"81ff06d4",
  1038 => x"0c535380",
  1039 => x"c7fc0885",
  1040 => x"3871892b",
  1041 => x"5271982a",
  1042 => x"d40c7190",
  1043 => x"2a7081ff",
  1044 => x"06d40c51",
  1045 => x"71882a70",
  1046 => x"81ff06d4",
  1047 => x"0c517181",
  1048 => x"ff06d40c",
  1049 => x"72902a70",
  1050 => x"81ff06d4",
  1051 => x"0c51d408",
  1052 => x"7081ff06",
  1053 => x"515182b8",
  1054 => x"bf527081",
  1055 => x"ff2e0981",
  1056 => x"06943881",
  1057 => x"ff0bd40c",
  1058 => x"d4087081",
  1059 => x"ff06ff14",
  1060 => x"54515171",
  1061 => x"e53870be",
  1062 => x"880c028c",
  1063 => x"050d0402",
  1064 => x"fc050d81",
  1065 => x"c75181ff",
  1066 => x"0bd40cff",
  1067 => x"11517080",
  1068 => x"25f43802",
  1069 => x"84050d04",
  1070 => x"02f0050d",
  1071 => x"a19f2d8f",
  1072 => x"cf538052",
  1073 => x"87fc80f7",
  1074 => x"51a0ad2d",
  1075 => x"be880854",
  1076 => x"be880881",
  1077 => x"2e098106",
  1078 => x"a33881ff",
  1079 => x"0bd40c82",
  1080 => x"0a52849c",
  1081 => x"80e951a0",
  1082 => x"ad2dbe88",
  1083 => x"088b3881",
  1084 => x"ff0bd40c",
  1085 => x"7353a282",
  1086 => x"04a19f2d",
  1087 => x"ff135372",
  1088 => x"c13872be",
  1089 => x"880c0290",
  1090 => x"050d0402",
  1091 => x"f4050d81",
  1092 => x"ff0bd40c",
  1093 => x"93538052",
  1094 => x"87fc80c1",
  1095 => x"51a0ad2d",
  1096 => x"be88088b",
  1097 => x"3881ff0b",
  1098 => x"d40c8153",
  1099 => x"a2b804a1",
  1100 => x"9f2dff13",
  1101 => x"5372df38",
  1102 => x"72be880c",
  1103 => x"028c050d",
  1104 => x"0402f005",
  1105 => x"0da19f2d",
  1106 => x"83aa5284",
  1107 => x"9c80c851",
  1108 => x"a0ad2dbe",
  1109 => x"8808812e",
  1110 => x"09810692",
  1111 => x"389fdf2d",
  1112 => x"be880883",
  1113 => x"ffff0653",
  1114 => x"7283aa2e",
  1115 => x"9738a28b",
  1116 => x"2da2ff04",
  1117 => x"8154a3e4",
  1118 => x"04ba9451",
  1119 => x"85f22d80",
  1120 => x"54a3e404",
  1121 => x"81ff0bd4",
  1122 => x"0cb153a1",
  1123 => x"b82dbe88",
  1124 => x"08802e80",
  1125 => x"c0388052",
  1126 => x"87fc80fa",
  1127 => x"51a0ad2d",
  1128 => x"be8808b1",
  1129 => x"3881ff0b",
  1130 => x"d40cd408",
  1131 => x"5381ff0b",
  1132 => x"d40c81ff",
  1133 => x"0bd40c81",
  1134 => x"ff0bd40c",
  1135 => x"81ff0bd4",
  1136 => x"0c72862a",
  1137 => x"708106be",
  1138 => x"88085651",
  1139 => x"5372802e",
  1140 => x"9338a2f4",
  1141 => x"0472822e",
  1142 => x"ff9f38ff",
  1143 => x"135372ff",
  1144 => x"aa387254",
  1145 => x"73be880c",
  1146 => x"0290050d",
  1147 => x"0402f005",
  1148 => x"0d810b80",
  1149 => x"c7fc0c84",
  1150 => x"54d00870",
  1151 => x"8f2a7081",
  1152 => x"06515153",
  1153 => x"72f33872",
  1154 => x"d00ca19f",
  1155 => x"2dbaa451",
  1156 => x"85f22dd0",
  1157 => x"08708f2a",
  1158 => x"70810651",
  1159 => x"515372f3",
  1160 => x"38810bd0",
  1161 => x"0cb15380",
  1162 => x"5284d480",
  1163 => x"c051a0ad",
  1164 => x"2dbe8808",
  1165 => x"812ea138",
  1166 => x"72822e09",
  1167 => x"81068c38",
  1168 => x"bab05185",
  1169 => x"f22d8053",
  1170 => x"a58e04ff",
  1171 => x"135372d7",
  1172 => x"38ff1454",
  1173 => x"73ffa238",
  1174 => x"a2c12dbe",
  1175 => x"880880c7",
  1176 => x"fc0cbe88",
  1177 => x"088b3881",
  1178 => x"5287fc80",
  1179 => x"d051a0ad",
  1180 => x"2d81ff0b",
  1181 => x"d40cd008",
  1182 => x"708f2a70",
  1183 => x"81065151",
  1184 => x"5372f338",
  1185 => x"72d00c81",
  1186 => x"ff0bd40c",
  1187 => x"815372be",
  1188 => x"880c0290",
  1189 => x"050d0402",
  1190 => x"e8050d78",
  1191 => x"5681ff0b",
  1192 => x"d40cd008",
  1193 => x"708f2a70",
  1194 => x"81065151",
  1195 => x"5372f338",
  1196 => x"82810bd0",
  1197 => x"0c81ff0b",
  1198 => x"d40c7752",
  1199 => x"87fc80d8",
  1200 => x"51a0ad2d",
  1201 => x"be880880",
  1202 => x"2e8c38ba",
  1203 => x"c85185f2",
  1204 => x"2d8153a6",
  1205 => x"ce0481ff",
  1206 => x"0bd40c81",
  1207 => x"fe0bd40c",
  1208 => x"80ff5575",
  1209 => x"70840557",
  1210 => x"0870982a",
  1211 => x"d40c7090",
  1212 => x"2c7081ff",
  1213 => x"06d40c54",
  1214 => x"70882c70",
  1215 => x"81ff06d4",
  1216 => x"0c547081",
  1217 => x"ff06d40c",
  1218 => x"54ff1555",
  1219 => x"748025d3",
  1220 => x"3881ff0b",
  1221 => x"d40c81ff",
  1222 => x"0bd40c81",
  1223 => x"ff0bd40c",
  1224 => x"868da054",
  1225 => x"81ff0bd4",
  1226 => x"0cd40881",
  1227 => x"ff065574",
  1228 => x"8738ff14",
  1229 => x"5473ed38",
  1230 => x"81ff0bd4",
  1231 => x"0cd00870",
  1232 => x"8f2a7081",
  1233 => x"06515153",
  1234 => x"72f33872",
  1235 => x"d00c72be",
  1236 => x"880c0298",
  1237 => x"050d0402",
  1238 => x"e8050d78",
  1239 => x"55805681",
  1240 => x"ff0bd40c",
  1241 => x"d008708f",
  1242 => x"2a708106",
  1243 => x"51515372",
  1244 => x"f3388281",
  1245 => x"0bd00c81",
  1246 => x"ff0bd40c",
  1247 => x"775287fc",
  1248 => x"80d151a0",
  1249 => x"ad2d80db",
  1250 => x"c6df54be",
  1251 => x"8808802e",
  1252 => x"8a38bad8",
  1253 => x"5185f22d",
  1254 => x"a7ee0481",
  1255 => x"ff0bd40c",
  1256 => x"d4087081",
  1257 => x"ff065153",
  1258 => x"7281fe2e",
  1259 => x"0981069d",
  1260 => x"3880ff53",
  1261 => x"9fdf2dbe",
  1262 => x"88087570",
  1263 => x"8405570c",
  1264 => x"ff135372",
  1265 => x"8025ed38",
  1266 => x"8156a7d3",
  1267 => x"04ff1454",
  1268 => x"73c93881",
  1269 => x"ff0bd40c",
  1270 => x"81ff0bd4",
  1271 => x"0cd00870",
  1272 => x"8f2a7081",
  1273 => x"06515153",
  1274 => x"72f33872",
  1275 => x"d00c75be",
  1276 => x"880c0298",
  1277 => x"050d0402",
  1278 => x"f4050d74",
  1279 => x"70882a83",
  1280 => x"fe800670",
  1281 => x"72982a07",
  1282 => x"72882b87",
  1283 => x"fc808006",
  1284 => x"73982b81",
  1285 => x"f00a0671",
  1286 => x"730707be",
  1287 => x"880c5651",
  1288 => x"5351028c",
  1289 => x"050d0402",
  1290 => x"f8050d02",
  1291 => x"8e0580f5",
  1292 => x"2d74882b",
  1293 => x"077083ff",
  1294 => x"ff06be88",
  1295 => x"0c510288",
  1296 => x"050d0402",
  1297 => x"fc050d72",
  1298 => x"5180710c",
  1299 => x"800b8412",
  1300 => x"0c028405",
  1301 => x"0d0402f0",
  1302 => x"050d7570",
  1303 => x"08841208",
  1304 => x"535353ff",
  1305 => x"5471712e",
  1306 => x"a838ac9a",
  1307 => x"2d841308",
  1308 => x"70842914",
  1309 => x"88117008",
  1310 => x"7081ff06",
  1311 => x"84180881",
  1312 => x"11870684",
  1313 => x"1a0c5351",
  1314 => x"55515151",
  1315 => x"ac942d71",
  1316 => x"5473be88",
  1317 => x"0c029005",
  1318 => x"0d0402f8",
  1319 => x"050dac9a",
  1320 => x"2de00870",
  1321 => x"8b2a7081",
  1322 => x"06515252",
  1323 => x"70802ea1",
  1324 => x"3880c880",
  1325 => x"08708429",
  1326 => x"80c88805",
  1327 => x"7381ff06",
  1328 => x"710c5151",
  1329 => x"80c88008",
  1330 => x"81118706",
  1331 => x"80c8800c",
  1332 => x"51800b80",
  1333 => x"c8a80cac",
  1334 => x"8d2dac94",
  1335 => x"2d028805",
  1336 => x"0d0402fc",
  1337 => x"050dac9a",
  1338 => x"2d810b80",
  1339 => x"c8a80cac",
  1340 => x"942d80c8",
  1341 => x"a8085170",
  1342 => x"f9380284",
  1343 => x"050d0402",
  1344 => x"fc050d80",
  1345 => x"c88051a8",
  1346 => x"c32da99a",
  1347 => x"51ac892d",
  1348 => x"abb32d02",
  1349 => x"84050d04",
  1350 => x"02f4050d",
  1351 => x"ab9a04be",
  1352 => x"880881f0",
  1353 => x"2e098106",
  1354 => x"8938810b",
  1355 => x"bdfc0cab",
  1356 => x"9a04be88",
  1357 => x"0881e02e",
  1358 => x"09810689",
  1359 => x"38810bbe",
  1360 => x"800cab9a",
  1361 => x"04be8808",
  1362 => x"52be8008",
  1363 => x"802e8838",
  1364 => x"be880881",
  1365 => x"80055271",
  1366 => x"842c728f",
  1367 => x"065353bd",
  1368 => x"fc08802e",
  1369 => x"99387284",
  1370 => x"29bdbc05",
  1371 => x"72138171",
  1372 => x"2b700973",
  1373 => x"0806730c",
  1374 => x"515353ab",
  1375 => x"90047284",
  1376 => x"29bdbc05",
  1377 => x"72138371",
  1378 => x"2b720807",
  1379 => x"720c5353",
  1380 => x"800bbe80",
  1381 => x"0c800bbd",
  1382 => x"fc0c80c8",
  1383 => x"8051a8d6",
  1384 => x"2dbe8808",
  1385 => x"ff24fef7",
  1386 => x"38800bbe",
  1387 => x"880c028c",
  1388 => x"050d0402",
  1389 => x"f8050dbd",
  1390 => x"bc528f51",
  1391 => x"80727084",
  1392 => x"05540cff",
  1393 => x"11517080",
  1394 => x"25f23802",
  1395 => x"88050d04",
  1396 => x"02f0050d",
  1397 => x"7551ac9a",
  1398 => x"2d70822c",
  1399 => x"fc06bdbc",
  1400 => x"1172109e",
  1401 => x"06710870",
  1402 => x"722a7083",
  1403 => x"0682742b",
  1404 => x"70097406",
  1405 => x"760c5451",
  1406 => x"56575351",
  1407 => x"53ac942d",
  1408 => x"71be880c",
  1409 => x"0290050d",
  1410 => x"0471980c",
  1411 => x"04ffb008",
  1412 => x"be880c04",
  1413 => x"810bffb0",
  1414 => x"0c04800b",
  1415 => x"ffb00c04",
  1416 => x"02fc050d",
  1417 => x"810bbe84",
  1418 => x"0c815184",
  1419 => x"e62d0284",
  1420 => x"050d0402",
  1421 => x"fc050d80",
  1422 => x"0bbe840c",
  1423 => x"805184e6",
  1424 => x"2d028405",
  1425 => x"0d0402ec",
  1426 => x"050d7654",
  1427 => x"8052870b",
  1428 => x"881580f5",
  1429 => x"2d565374",
  1430 => x"72248338",
  1431 => x"a0537251",
  1432 => x"82ef2d81",
  1433 => x"128b1580",
  1434 => x"f52d5452",
  1435 => x"727225de",
  1436 => x"38029405",
  1437 => x"0d0402f0",
  1438 => x"050d80c8",
  1439 => x"b8085481",
  1440 => x"f82d800b",
  1441 => x"80c8bc0c",
  1442 => x"7308802e",
  1443 => x"81843882",
  1444 => x"0bbe9c0c",
  1445 => x"80c8bc08",
  1446 => x"8f06be98",
  1447 => x"0c730852",
  1448 => x"71832e96",
  1449 => x"38718326",
  1450 => x"89387181",
  1451 => x"2eaf38ad",
  1452 => x"fb047185",
  1453 => x"2e9f38ad",
  1454 => x"fb048814",
  1455 => x"80f52d84",
  1456 => x"1508bae8",
  1457 => x"53545285",
  1458 => x"f22d7184",
  1459 => x"29137008",
  1460 => x"5252adff",
  1461 => x"047351ac",
  1462 => x"c62dadfb",
  1463 => x"0480c8ac",
  1464 => x"08881508",
  1465 => x"2c708106",
  1466 => x"51527180",
  1467 => x"2e8738ba",
  1468 => x"ec51adf8",
  1469 => x"04baf051",
  1470 => x"85f22d84",
  1471 => x"14085185",
  1472 => x"f22d80c8",
  1473 => x"bc088105",
  1474 => x"80c8bc0c",
  1475 => x"8c1454ad",
  1476 => x"88040290",
  1477 => x"050d0471",
  1478 => x"80c8b80c",
  1479 => x"acf62d80",
  1480 => x"c8bc08ff",
  1481 => x"0580c8c0",
  1482 => x"0c047180",
  1483 => x"c8c40c04",
  1484 => x"02e8050d",
  1485 => x"80c8b808",
  1486 => x"80c8c408",
  1487 => x"575580f8",
  1488 => x"51abd02d",
  1489 => x"be880881",
  1490 => x"2a708106",
  1491 => x"5152719b",
  1492 => x"388751ab",
  1493 => x"d02dbe88",
  1494 => x"08812a70",
  1495 => x"81065152",
  1496 => x"71802eb1",
  1497 => x"38aeeb04",
  1498 => x"aa982d87",
  1499 => x"51abd02d",
  1500 => x"be8808f4",
  1501 => x"38aefb04",
  1502 => x"aa982d80",
  1503 => x"f851abd0",
  1504 => x"2dbe8808",
  1505 => x"f338be84",
  1506 => x"08813270",
  1507 => x"be840c70",
  1508 => x"525284e6",
  1509 => x"2d800b80",
  1510 => x"c8b00c80",
  1511 => x"0b80c8b4",
  1512 => x"0cbe8408",
  1513 => x"82fd3880",
  1514 => x"da51abd0",
  1515 => x"2dbe8808",
  1516 => x"802e8c38",
  1517 => x"80c8b008",
  1518 => x"81800780",
  1519 => x"c8b00c80",
  1520 => x"d951abd0",
  1521 => x"2dbe8808",
  1522 => x"802e8c38",
  1523 => x"80c8b008",
  1524 => x"80c00780",
  1525 => x"c8b00c81",
  1526 => x"9451abd0",
  1527 => x"2dbe8808",
  1528 => x"802e8b38",
  1529 => x"80c8b008",
  1530 => x"900780c8",
  1531 => x"b00c8191",
  1532 => x"51abd02d",
  1533 => x"be880880",
  1534 => x"2e8b3880",
  1535 => x"c8b008a0",
  1536 => x"0780c8b0",
  1537 => x"0c81f551",
  1538 => x"abd02dbe",
  1539 => x"8808802e",
  1540 => x"8b3880c8",
  1541 => x"b0088107",
  1542 => x"80c8b00c",
  1543 => x"81f251ab",
  1544 => x"d02dbe88",
  1545 => x"08802e8b",
  1546 => x"3880c8b0",
  1547 => x"08820780",
  1548 => x"c8b00c81",
  1549 => x"eb51abd0",
  1550 => x"2dbe8808",
  1551 => x"802e8b38",
  1552 => x"80c8b008",
  1553 => x"840780c8",
  1554 => x"b00c81f4",
  1555 => x"51abd02d",
  1556 => x"be880880",
  1557 => x"2e8b3880",
  1558 => x"c8b00888",
  1559 => x"0780c8b0",
  1560 => x"0c80d851",
  1561 => x"abd02dbe",
  1562 => x"8808802e",
  1563 => x"8c3880c8",
  1564 => x"b4088180",
  1565 => x"0780c8b4",
  1566 => x"0c9251ab",
  1567 => x"d02dbe88",
  1568 => x"08802e8c",
  1569 => x"3880c8b4",
  1570 => x"0880c007",
  1571 => x"80c8b40c",
  1572 => x"9451abd0",
  1573 => x"2dbe8808",
  1574 => x"802e8b38",
  1575 => x"80c8b408",
  1576 => x"900780c8",
  1577 => x"b40c9151",
  1578 => x"abd02dbe",
  1579 => x"8808802e",
  1580 => x"8b3880c8",
  1581 => x"b408a007",
  1582 => x"80c8b40c",
  1583 => x"9d51abd0",
  1584 => x"2dbe8808",
  1585 => x"802e8b38",
  1586 => x"80c8b408",
  1587 => x"810780c8",
  1588 => x"b40c9b51",
  1589 => x"abd02dbe",
  1590 => x"8808802e",
  1591 => x"8b3880c8",
  1592 => x"b4088207",
  1593 => x"80c8b40c",
  1594 => x"9c51abd0",
  1595 => x"2dbe8808",
  1596 => x"802e8b38",
  1597 => x"80c8b408",
  1598 => x"840780c8",
  1599 => x"b40ca351",
  1600 => x"abd02dbe",
  1601 => x"8808802e",
  1602 => x"8b3880c8",
  1603 => x"b4088807",
  1604 => x"80c8b40c",
  1605 => x"81fd51ab",
  1606 => x"d02d81fa",
  1607 => x"51abd02d",
  1608 => x"b7eb0481",
  1609 => x"f551abd0",
  1610 => x"2dbe8808",
  1611 => x"812a7081",
  1612 => x"06515271",
  1613 => x"802eb338",
  1614 => x"80c8c008",
  1615 => x"5271802e",
  1616 => x"8a38ff12",
  1617 => x"80c8c00c",
  1618 => x"b2ea0480",
  1619 => x"c8bc0810",
  1620 => x"80c8bc08",
  1621 => x"05708429",
  1622 => x"16515288",
  1623 => x"1208802e",
  1624 => x"8938ff51",
  1625 => x"88120852",
  1626 => x"712d81f2",
  1627 => x"51abd02d",
  1628 => x"be880881",
  1629 => x"2a708106",
  1630 => x"51527180",
  1631 => x"2eb43880",
  1632 => x"c8bc08ff",
  1633 => x"1180c8c0",
  1634 => x"08565353",
  1635 => x"7372258a",
  1636 => x"38811480",
  1637 => x"c8c00cb3",
  1638 => x"b2047210",
  1639 => x"13708429",
  1640 => x"16515288",
  1641 => x"1208802e",
  1642 => x"8938fe51",
  1643 => x"88120852",
  1644 => x"712d81fd",
  1645 => x"51abd02d",
  1646 => x"be880881",
  1647 => x"2a708106",
  1648 => x"51527180",
  1649 => x"2eb13880",
  1650 => x"c8c00880",
  1651 => x"2e8a3880",
  1652 => x"0b80c8c0",
  1653 => x"0cb3f704",
  1654 => x"80c8bc08",
  1655 => x"1080c8bc",
  1656 => x"08057084",
  1657 => x"29165152",
  1658 => x"88120880",
  1659 => x"2e8938fd",
  1660 => x"51881208",
  1661 => x"52712d81",
  1662 => x"fa51abd0",
  1663 => x"2dbe8808",
  1664 => x"812a7081",
  1665 => x"06515271",
  1666 => x"802eb138",
  1667 => x"80c8bc08",
  1668 => x"ff115452",
  1669 => x"80c8c008",
  1670 => x"73258938",
  1671 => x"7280c8c0",
  1672 => x"0cb4bc04",
  1673 => x"71101270",
  1674 => x"84291651",
  1675 => x"52881208",
  1676 => x"802e8938",
  1677 => x"fc518812",
  1678 => x"0852712d",
  1679 => x"80c8c008",
  1680 => x"70535473",
  1681 => x"802e8a38",
  1682 => x"8c15ff15",
  1683 => x"5555b4c3",
  1684 => x"04820bbe",
  1685 => x"9c0c718f",
  1686 => x"06be980c",
  1687 => x"81eb51ab",
  1688 => x"d02dbe88",
  1689 => x"08812a70",
  1690 => x"81065152",
  1691 => x"71802ead",
  1692 => x"38740885",
  1693 => x"2e098106",
  1694 => x"a4388815",
  1695 => x"80f52dff",
  1696 => x"05527188",
  1697 => x"1681b72d",
  1698 => x"71982b52",
  1699 => x"71802588",
  1700 => x"38800b88",
  1701 => x"1681b72d",
  1702 => x"7451acc6",
  1703 => x"2d81f451",
  1704 => x"abd02dbe",
  1705 => x"8808812a",
  1706 => x"70810651",
  1707 => x"5271802e",
  1708 => x"b3387408",
  1709 => x"852e0981",
  1710 => x"06aa3888",
  1711 => x"1580f52d",
  1712 => x"81055271",
  1713 => x"881681b7",
  1714 => x"2d7181ff",
  1715 => x"068b1680",
  1716 => x"f52d5452",
  1717 => x"72722787",
  1718 => x"38728816",
  1719 => x"81b72d74",
  1720 => x"51acc62d",
  1721 => x"80da51ab",
  1722 => x"d02dbe88",
  1723 => x"08812a70",
  1724 => x"81065152",
  1725 => x"71802e81",
  1726 => x"ac3880c8",
  1727 => x"b80880c8",
  1728 => x"c0085553",
  1729 => x"73802e8a",
  1730 => x"388c13ff",
  1731 => x"155553b6",
  1732 => x"84047208",
  1733 => x"5271822e",
  1734 => x"a6387182",
  1735 => x"26893871",
  1736 => x"812eaa38",
  1737 => x"b7a50471",
  1738 => x"832eb438",
  1739 => x"71842e09",
  1740 => x"810680f1",
  1741 => x"38881308",
  1742 => x"51ae972d",
  1743 => x"b7a50480",
  1744 => x"c8c00851",
  1745 => x"88130852",
  1746 => x"712db7a5",
  1747 => x"04810b88",
  1748 => x"14082b80",
  1749 => x"c8ac0832",
  1750 => x"80c8ac0c",
  1751 => x"b6fa0488",
  1752 => x"1380f52d",
  1753 => x"81058b14",
  1754 => x"80f52d53",
  1755 => x"54717424",
  1756 => x"83388054",
  1757 => x"73881481",
  1758 => x"b72dacf6",
  1759 => x"2db7a504",
  1760 => x"7508802e",
  1761 => x"a3387508",
  1762 => x"51abd02d",
  1763 => x"be880881",
  1764 => x"06527180",
  1765 => x"2e8c3880",
  1766 => x"c8c00851",
  1767 => x"84160852",
  1768 => x"712d8816",
  1769 => x"5675d938",
  1770 => x"8054800b",
  1771 => x"be9c0c73",
  1772 => x"8f06be98",
  1773 => x"0ca05273",
  1774 => x"80c8c008",
  1775 => x"2e098106",
  1776 => x"993880c8",
  1777 => x"bc08ff05",
  1778 => x"74327009",
  1779 => x"81057072",
  1780 => x"079f2a91",
  1781 => x"71315151",
  1782 => x"53537151",
  1783 => x"82ef2d81",
  1784 => x"14548e74",
  1785 => x"25c438be",
  1786 => x"84085271",
  1787 => x"be880c02",
  1788 => x"98050d04",
  1789 => x"00ffffff",
  1790 => x"ff00ffff",
  1791 => x"ffff00ff",
  1792 => x"ffffff00",
  1793 => x"52657365",
  1794 => x"74000000",
  1795 => x"53617665",
  1796 => x"20736574",
  1797 => x"74696e67",
  1798 => x"73000000",
  1799 => x"5363616e",
  1800 => x"6c696e65",
  1801 => x"73000000",
  1802 => x"4c6f6164",
  1803 => x"20524f4d",
  1804 => x"20100000",
  1805 => x"45786974",
  1806 => x"00000000",
  1807 => x"50432045",
  1808 => x"6e67696e",
  1809 => x"65206d6f",
  1810 => x"64650000",
  1811 => x"54757262",
  1812 => x"6f677261",
  1813 => x"66782031",
  1814 => x"36206d6f",
  1815 => x"64650000",
  1816 => x"56474120",
  1817 => x"2d203331",
  1818 => x"4b487a2c",
  1819 => x"20363048",
  1820 => x"7a000000",
  1821 => x"5456202d",
  1822 => x"20343830",
  1823 => x"692c2036",
  1824 => x"30487a00",
  1825 => x"4261636b",
  1826 => x"00000000",
  1827 => x"46504741",
  1828 => x"50434520",
  1829 => x"43464700",
  1830 => x"496e6974",
  1831 => x"69616c69",
  1832 => x"7a696e67",
  1833 => x"20534420",
  1834 => x"63617264",
  1835 => x"0a000000",
  1836 => x"424f4f54",
  1837 => x"20202020",
  1838 => x"50434500",
  1839 => x"43617264",
  1840 => x"20696e69",
  1841 => x"74206661",
  1842 => x"696c6564",
  1843 => x"0a000000",
  1844 => x"4d425220",
  1845 => x"6661696c",
  1846 => x"0a000000",
  1847 => x"46415431",
  1848 => x"36202020",
  1849 => x"00000000",
  1850 => x"46415433",
  1851 => x"32202020",
  1852 => x"00000000",
  1853 => x"4e6f2070",
  1854 => x"61727469",
  1855 => x"74696f6e",
  1856 => x"20736967",
  1857 => x"0a000000",
  1858 => x"42616420",
  1859 => x"70617274",
  1860 => x"0a000000",
  1861 => x"53444843",
  1862 => x"20657272",
  1863 => x"6f72210a",
  1864 => x"00000000",
  1865 => x"53442069",
  1866 => x"6e69742e",
  1867 => x"2e2e0a00",
  1868 => x"53442063",
  1869 => x"61726420",
  1870 => x"72657365",
  1871 => x"74206661",
  1872 => x"696c6564",
  1873 => x"210a0000",
  1874 => x"57726974",
  1875 => x"65206661",
  1876 => x"696c6564",
  1877 => x"0a000000",
  1878 => x"52656164",
  1879 => x"20666169",
  1880 => x"6c65640a",
  1881 => x"00000000",
  1882 => x"16200000",
  1883 => x"14200000",
  1884 => x"15200000",
  1885 => x"00000002",
  1886 => x"00000002",
  1887 => x"00001c04",
  1888 => x"000004c0",
  1889 => x"00000002",
  1890 => x"00001c0c",
  1891 => x"0000037d",
  1892 => x"00000003",
  1893 => x"00001de0",
  1894 => x"00000002",
  1895 => x"00000001",
  1896 => x"00001c1c",
  1897 => x"00000001",
  1898 => x"00000003",
  1899 => x"00001dd8",
  1900 => x"00000002",
  1901 => x"00000002",
  1902 => x"00001c28",
  1903 => x"00000786",
  1904 => x"00000002",
  1905 => x"00001c34",
  1906 => x"00001633",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00001c3c",
  1911 => x"00001c4c",
  1912 => x"00001c60",
  1913 => x"00001c74",
  1914 => x"0000004d",
  1915 => x"0000075a",
  1916 => x"0000002c",
  1917 => x"00000770",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000002",
  1921 => x"00001f38",
  1922 => x"0000054e",
  1923 => x"00000002",
  1924 => x"00001f56",
  1925 => x"0000054e",
  1926 => x"00000002",
  1927 => x"00001f74",
  1928 => x"0000054e",
  1929 => x"00000002",
  1930 => x"00001f92",
  1931 => x"0000054e",
  1932 => x"00000002",
  1933 => x"00001fb0",
  1934 => x"0000054e",
  1935 => x"00000002",
  1936 => x"00001fce",
  1937 => x"0000054e",
  1938 => x"00000002",
  1939 => x"00001fec",
  1940 => x"0000054e",
  1941 => x"00000002",
  1942 => x"0000200a",
  1943 => x"0000054e",
  1944 => x"00000002",
  1945 => x"00002028",
  1946 => x"0000054e",
  1947 => x"00000002",
  1948 => x"00002046",
  1949 => x"0000054e",
  1950 => x"00000002",
  1951 => x"00002064",
  1952 => x"0000054e",
  1953 => x"00000002",
  1954 => x"00002082",
  1955 => x"0000054e",
  1956 => x"00000002",
  1957 => x"000020a0",
  1958 => x"0000054e",
  1959 => x"00000004",
  1960 => x"00001c84",
  1961 => x"00001d78",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"000006ee",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

