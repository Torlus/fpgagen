-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"000b0b0b",
     4 => x"0b8c04ff",
     5 => x"0d800404",
     6 => x"00000017",
     7 => x"00000000",
     8 => x"0b0b80c0",
     9 => x"e4080b0b",
    10 => x"80c0e808",
    11 => x"0b0b80c0",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c0ec0c0b",
    16 => x"0b80c0e8",
    17 => x"0c0b0b80",
    18 => x"c0e40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bba98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c0e470",
    57 => x"80cba427",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c519098",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c0",
    65 => x"f40c9f0b",
    66 => x"80c0f80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c0f808ff",
    70 => x"0580c0f8",
    71 => x"0c80c0f8",
    72 => x"088025e8",
    73 => x"3880c0f4",
    74 => x"08ff0580",
    75 => x"c0f40c80",
    76 => x"c0f40880",
    77 => x"25d03802",
    78 => x"84050d04",
    79 => x"02f0050d",
    80 => x"f88053f8",
    81 => x"a05483bf",
    82 => x"52737081",
    83 => x"05553351",
    84 => x"70737081",
    85 => x"055534ff",
    86 => x"12527180",
    87 => x"25eb38fb",
    88 => x"c0539f52",
    89 => x"a0737081",
    90 => x"055534ff",
    91 => x"12527180",
    92 => x"25f23802",
    93 => x"90050d04",
    94 => x"02f4050d",
    95 => x"74538e0b",
    96 => x"80c0f408",
    97 => x"25913882",
    98 => x"bc2d80c0",
    99 => x"f408ff05",
   100 => x"80c0f40c",
   101 => x"82fe0480",
   102 => x"c0f40880",
   103 => x"c0f80853",
   104 => x"51728a2e",
   105 => x"098106be",
   106 => x"38715171",
   107 => x"9f24a438",
   108 => x"80c0f408",
   109 => x"a02911f8",
   110 => x"80115151",
   111 => x"a0713480",
   112 => x"c0f80881",
   113 => x"0580c0f8",
   114 => x"0c80c0f8",
   115 => x"08519f71",
   116 => x"25de3880",
   117 => x"0b80c0f8",
   118 => x"0c80c0f4",
   119 => x"08810580",
   120 => x"c0f40c83",
   121 => x"fc0470a0",
   122 => x"2912f880",
   123 => x"11515172",
   124 => x"713480c0",
   125 => x"f8088105",
   126 => x"80c0f80c",
   127 => x"80c0f808",
   128 => x"a02e0981",
   129 => x"06913880",
   130 => x"0b80c0f8",
   131 => x"0c80c0f4",
   132 => x"08810580",
   133 => x"c0f40c02",
   134 => x"8c050d04",
   135 => x"02e8050d",
   136 => x"77795656",
   137 => x"880bfc16",
   138 => x"77712c8f",
   139 => x"06545254",
   140 => x"80537272",
   141 => x"25953871",
   142 => x"53fbe014",
   143 => x"51877134",
   144 => x"8114ff14",
   145 => x"545472f1",
   146 => x"387153f9",
   147 => x"1576712c",
   148 => x"87065351",
   149 => x"71802e8b",
   150 => x"38fbe014",
   151 => x"51717134",
   152 => x"81145472",
   153 => x"8e249538",
   154 => x"8f733153",
   155 => x"fbe01451",
   156 => x"a0713481",
   157 => x"14ff1454",
   158 => x"5472f138",
   159 => x"0298050d",
   160 => x"0402ec05",
   161 => x"0d800b80",
   162 => x"c0fc0cf6",
   163 => x"8c08f690",
   164 => x"0871882c",
   165 => x"565481ff",
   166 => x"06527372",
   167 => x"25893871",
   168 => x"54820b80",
   169 => x"c0fc0c72",
   170 => x"882c7381",
   171 => x"ff065455",
   172 => x"7473258d",
   173 => x"387280c0",
   174 => x"fc088407",
   175 => x"80c0fc0c",
   176 => x"5573842b",
   177 => x"87e87125",
   178 => x"83713170",
   179 => x"0b0b0bbd",
   180 => x"a80c8171",
   181 => x"2bf6880c",
   182 => x"fea413ff",
   183 => x"122c7888",
   184 => x"29ff9405",
   185 => x"70812c80",
   186 => x"c0fc0852",
   187 => x"58525551",
   188 => x"52547680",
   189 => x"2e853870",
   190 => x"81075170",
   191 => x"f6940c71",
   192 => x"098105f6",
   193 => x"800c7209",
   194 => x"8105f684",
   195 => x"0c029405",
   196 => x"0d0402f4",
   197 => x"050d7453",
   198 => x"72708105",
   199 => x"5480f52d",
   200 => x"5271802e",
   201 => x"89387151",
   202 => x"82f82d86",
   203 => x"9804028c",
   204 => x"050d0402",
   205 => x"f4050d74",
   206 => x"70820680",
   207 => x"cb880cbd",
   208 => x"c8718106",
   209 => x"54545171",
   210 => x"881481b7",
   211 => x"2d70822a",
   212 => x"70810651",
   213 => x"5170a014",
   214 => x"81b72d70",
   215 => x"80c0e40c",
   216 => x"028c050d",
   217 => x"0402f805",
   218 => x"0dbbc052",
   219 => x"80c18051",
   220 => x"9e932d80",
   221 => x"c0e40880",
   222 => x"2ea33880",
   223 => x"c49c5280",
   224 => x"c18051a0",
   225 => x"e02d80c4",
   226 => x"9c0880c1",
   227 => x"8c0c80c4",
   228 => x"9c08fec0",
   229 => x"0c80c49c",
   230 => x"085186b3",
   231 => x"2d028805",
   232 => x"0d0402f0",
   233 => x"050d8051",
   234 => x"93c72dbb",
   235 => x"c05280c1",
   236 => x"80519e93",
   237 => x"2d80c0e4",
   238 => x"08802eaa",
   239 => x"3880c18c",
   240 => x"0880c49c",
   241 => x"0c80c4a0",
   242 => x"5480fd53",
   243 => x"80747084",
   244 => x"05560cff",
   245 => x"13537280",
   246 => x"25f23880",
   247 => x"c49c5280",
   248 => x"c18051a1",
   249 => x"892d0290",
   250 => x"050d0402",
   251 => x"d8050d80",
   252 => x"0bbdac0c",
   253 => x"80c18c08",
   254 => x"fec00c81",
   255 => x"0bfec40c",
   256 => x"840bfec4",
   257 => x"0c7b5280",
   258 => x"c180519e",
   259 => x"932d80c0",
   260 => x"e4085380",
   261 => x"c0e40880",
   262 => x"2e81b838",
   263 => x"80c18408",
   264 => x"55800bff",
   265 => x"16575975",
   266 => x"792e8b38",
   267 => x"81197681",
   268 => x"2a575975",
   269 => x"f738f719",
   270 => x"5974b080",
   271 => x"802e0981",
   272 => x"06893882",
   273 => x"0bfedc0c",
   274 => x"88e20474",
   275 => x"9880802e",
   276 => x"09810689",
   277 => x"38810bfe",
   278 => x"dc0c88e2",
   279 => x"04800bfe",
   280 => x"dc0c815a",
   281 => x"80752580",
   282 => x"e3387852",
   283 => x"7551849c",
   284 => x"2d80c49c",
   285 => x"5280c180",
   286 => x"51a0e02d",
   287 => x"80c0e408",
   288 => x"802ea838",
   289 => x"80c49c58",
   290 => x"83fc5777",
   291 => x"70840559",
   292 => x"087083ff",
   293 => x"ff067190",
   294 => x"2afec80c",
   295 => x"fec80cfc",
   296 => x"18585376",
   297 => x"8025e438",
   298 => x"89b30480",
   299 => x"c0e4085a",
   300 => x"84805580",
   301 => x"c18051a0",
   302 => x"b02dfc80",
   303 => x"15811757",
   304 => x"55748024",
   305 => x"ffa43879",
   306 => x"802e8638",
   307 => x"820bbdac",
   308 => x"0c795372",
   309 => x"80c0e40c",
   310 => x"02a8050d",
   311 => x"0402fc05",
   312 => x"0daeb42d",
   313 => x"fec45181",
   314 => x"710c8271",
   315 => x"0c028405",
   316 => x"0d0402f4",
   317 => x"050d7476",
   318 => x"78535452",
   319 => x"80712597",
   320 => x"38727081",
   321 => x"055480f5",
   322 => x"2d727081",
   323 => x"055481b7",
   324 => x"2dff1151",
   325 => x"70eb3880",
   326 => x"7281b72d",
   327 => x"028c050d",
   328 => x"0402e805",
   329 => x"0d775680",
   330 => x"70565473",
   331 => x"7624b638",
   332 => x"80caac08",
   333 => x"742eae38",
   334 => x"73519bd8",
   335 => x"2d80c0e4",
   336 => x"0880c0e4",
   337 => x"08098105",
   338 => x"7080c0e4",
   339 => x"08079f2a",
   340 => x"77058117",
   341 => x"57575353",
   342 => x"74762489",
   343 => x"3880caac",
   344 => x"087426d4",
   345 => x"387280c0",
   346 => x"e40c0298",
   347 => x"050d0402",
   348 => x"f4050dbf",
   349 => x"e0081551",
   350 => x"8aa12d80",
   351 => x"c0e40880",
   352 => x"2eac388b",
   353 => x"5380c0e4",
   354 => x"085280c8",
   355 => x"9c5189f2",
   356 => x"2d80c89c",
   357 => x"5187eb2d",
   358 => x"80c0e408",
   359 => x"802e8f38",
   360 => x"bdb051b0",
   361 => x"9b2daeb4",
   362 => x"2d80518b",
   363 => x"b904bfe4",
   364 => x"51b09b2d",
   365 => x"aea02d81",
   366 => x"5185812d",
   367 => x"028c050d",
   368 => x"0402dc05",
   369 => x"0d80705a",
   370 => x"5574bfe0",
   371 => x"0825b338",
   372 => x"80caac08",
   373 => x"752eab38",
   374 => x"78519bd8",
   375 => x"2d80c0e4",
   376 => x"08098105",
   377 => x"7080c0e4",
   378 => x"08079f2a",
   379 => x"7605811b",
   380 => x"5b565474",
   381 => x"bfe00825",
   382 => x"893880ca",
   383 => x"ac087926",
   384 => x"d7388055",
   385 => x"7880caac",
   386 => x"082781d9",
   387 => x"3878519b",
   388 => x"d82d80c0",
   389 => x"e408802e",
   390 => x"81ab3880",
   391 => x"c0e4088b",
   392 => x"0580f52d",
   393 => x"70842a70",
   394 => x"81067710",
   395 => x"78842b80",
   396 => x"c89c0b80",
   397 => x"f52d5c5c",
   398 => x"53515556",
   399 => x"73802e80",
   400 => x"ca387416",
   401 => x"822b8e89",
   402 => x"0bbeb412",
   403 => x"0c547775",
   404 => x"311080c1",
   405 => x"94115556",
   406 => x"90747081",
   407 => x"055681b7",
   408 => x"2da07481",
   409 => x"b72d7681",
   410 => x"ff068116",
   411 => x"58547380",
   412 => x"2e8a389c",
   413 => x"5380c89c",
   414 => x"528d8304",
   415 => x"8b5380c0",
   416 => x"e4085280",
   417 => x"c1961651",
   418 => x"8dbd0474",
   419 => x"16822b8a",
   420 => x"ef0bbeb4",
   421 => x"120c5476",
   422 => x"81ff0681",
   423 => x"16585473",
   424 => x"802e8a38",
   425 => x"9c5380c8",
   426 => x"9c528db4",
   427 => x"048b5380",
   428 => x"c0e40852",
   429 => x"77753110",
   430 => x"80c19405",
   431 => x"51765589",
   432 => x"f22d8dda",
   433 => x"04749029",
   434 => x"75317010",
   435 => x"80c19405",
   436 => x"515480c0",
   437 => x"e4087481",
   438 => x"b72d8119",
   439 => x"59748b24",
   440 => x"a3388c84",
   441 => x"04749029",
   442 => x"75317010",
   443 => x"80c19405",
   444 => x"8c773157",
   445 => x"51548074",
   446 => x"81b72d9e",
   447 => x"14ff1656",
   448 => x"5474f338",
   449 => x"02a4050d",
   450 => x"0402fc05",
   451 => x"0dbfe008",
   452 => x"13518aa1",
   453 => x"2d80c0e4",
   454 => x"08802e89",
   455 => x"3880c0e4",
   456 => x"085193c7",
   457 => x"2d800bbf",
   458 => x"e00c8bc1",
   459 => x"2daef82d",
   460 => x"0284050d",
   461 => x"0402fc05",
   462 => x"0d725170",
   463 => x"fd2ead38",
   464 => x"70fd248a",
   465 => x"3870fc2e",
   466 => x"80c4388f",
   467 => x"960470fe",
   468 => x"2eb13870",
   469 => x"ff2e0981",
   470 => x"06bc38bf",
   471 => x"e0085170",
   472 => x"802eb338",
   473 => x"ff11bfe0",
   474 => x"0c8f9604",
   475 => x"bfe008f0",
   476 => x"0570bfe0",
   477 => x"0c517080",
   478 => x"259c3880",
   479 => x"0bbfe00c",
   480 => x"8f9604bf",
   481 => x"e0088105",
   482 => x"bfe00c8f",
   483 => x"9604bfe0",
   484 => x"089005bf",
   485 => x"e00c8bc1",
   486 => x"2daef82d",
   487 => x"0284050d",
   488 => x"0402fc05",
   489 => x"0d800bbf",
   490 => x"e00c8bc1",
   491 => x"2dbeac51",
   492 => x"b09b2d02",
   493 => x"84050d04",
   494 => x"bdf40b80",
   495 => x"f52d80c0",
   496 => x"e40c0402",
   497 => x"fc050d72",
   498 => x"87065170",
   499 => x"bdf40b81",
   500 => x"b72d0284",
   501 => x"050d0402",
   502 => x"f8050d80",
   503 => x"cb880882",
   504 => x"06bdd00b",
   505 => x"80f52d52",
   506 => x"5270802e",
   507 => x"85387181",
   508 => x"0752bde8",
   509 => x"0b80f52d",
   510 => x"5170802e",
   511 => x"85387184",
   512 => x"075280c1",
   513 => x"9008802e",
   514 => x"85387190",
   515 => x"07527180",
   516 => x"c0e40c02",
   517 => x"88050d04",
   518 => x"02f0050d",
   519 => x"810b80c1",
   520 => x"900c800b",
   521 => x"bdac0c87",
   522 => x"53905186",
   523 => x"b32d7251",
   524 => x"8fc32d81",
   525 => x"0bfec40c",
   526 => x"840bfec4",
   527 => x"0c830bfe",
   528 => x"cc0cbbcc",
   529 => x"5186922d",
   530 => x"8452a5cf",
   531 => x"2d94ed2d",
   532 => x"80c0e408",
   533 => x"802e8638",
   534 => x"fe5290e5",
   535 => x"04ff1252",
   536 => x"718024e6",
   537 => x"3871802e",
   538 => x"828d38ab",
   539 => x"ed2dae94",
   540 => x"2dabd02d",
   541 => x"abd02d81",
   542 => x"f92d8151",
   543 => x"85812dab",
   544 => x"d02dabd0",
   545 => x"2d815185",
   546 => x"812d86e5",
   547 => x"2dbbe451",
   548 => x"87eb2d80",
   549 => x"c0e40880",
   550 => x"2e9438bd",
   551 => x"b051b09b",
   552 => x"2d805185",
   553 => x"812d820b",
   554 => x"bdac0c91",
   555 => x"b90480c0",
   556 => x"e408518f",
   557 => x"a12daea0",
   558 => x"2dac862d",
   559 => x"b0ae2d80",
   560 => x"c0e40880",
   561 => x"cb8c0888",
   562 => x"2b80cb90",
   563 => x"0807fed8",
   564 => x"0c548fd7",
   565 => x"2d80c0e4",
   566 => x"0880c18c",
   567 => x"082ea538",
   568 => x"80c0e408",
   569 => x"80c18c0c",
   570 => x"80c0e408",
   571 => x"fec00c84",
   572 => x"52735185",
   573 => x"812dabd0",
   574 => x"2dabd02d",
   575 => x"ff125271",
   576 => x"8025ee38",
   577 => x"8551adcd",
   578 => x"2d80c0e4",
   579 => x"08812a70",
   580 => x"81065152",
   581 => x"71802e95",
   582 => x"38ff1370",
   583 => x"09709f2c",
   584 => x"72067054",
   585 => x"5253538f",
   586 => x"c32daef8",
   587 => x"2d8651ad",
   588 => x"cd2d80c0",
   589 => x"e408812a",
   590 => x"70810651",
   591 => x"5271802e",
   592 => x"93388113",
   593 => x"53877325",
   594 => x"83388753",
   595 => x"72518fc3",
   596 => x"2daef82d",
   597 => x"8fb82d80",
   598 => x"c0e408fe",
   599 => x"d40c7380",
   600 => x"2e8c38bd",
   601 => x"ac088807",
   602 => x"fec40c91",
   603 => x"b904bdac",
   604 => x"08fec40c",
   605 => x"91b904bb",
   606 => x"f0518692",
   607 => x"2d800b80",
   608 => x"c0e40c02",
   609 => x"90050d04",
   610 => x"02e8050d",
   611 => x"77797b58",
   612 => x"55558053",
   613 => x"727625a3",
   614 => x"38747081",
   615 => x"055680f5",
   616 => x"2d747081",
   617 => x"055680f5",
   618 => x"2d525271",
   619 => x"712e8638",
   620 => x"815193bd",
   621 => x"04811353",
   622 => x"93940480",
   623 => x"517080c0",
   624 => x"e40c0298",
   625 => x"050d0402",
   626 => x"ec050d76",
   627 => x"5574802e",
   628 => x"80c2389a",
   629 => x"1580e02d",
   630 => x"51aa932d",
   631 => x"80c0e408",
   632 => x"80c0e408",
   633 => x"80cacc0c",
   634 => x"80c0e408",
   635 => x"545480ca",
   636 => x"a808802e",
   637 => x"9a389415",
   638 => x"80e02d51",
   639 => x"aa932d80",
   640 => x"c0e40890",
   641 => x"2b83fff0",
   642 => x"0a067075",
   643 => x"07515372",
   644 => x"80cacc0c",
   645 => x"80cacc08",
   646 => x"5372802e",
   647 => x"9d3880ca",
   648 => x"a008fe14",
   649 => x"712980ca",
   650 => x"b4080580",
   651 => x"cad00c70",
   652 => x"842b80ca",
   653 => x"ac0c5494",
   654 => x"e80480ca",
   655 => x"b80880ca",
   656 => x"cc0c80ca",
   657 => x"bc0880ca",
   658 => x"d00c80ca",
   659 => x"a808802e",
   660 => x"8b3880ca",
   661 => x"a008842b",
   662 => x"5394e304",
   663 => x"80cac008",
   664 => x"842b5372",
   665 => x"80caac0c",
   666 => x"0294050d",
   667 => x"0402d805",
   668 => x"0d800b80",
   669 => x"caa80c80",
   670 => x"c49c5280",
   671 => x"51a8bf2d",
   672 => x"80c0e408",
   673 => x"5480c0e4",
   674 => x"088c38bc",
   675 => x"84518692",
   676 => x"2d73559a",
   677 => x"d5048056",
   678 => x"810b80ca",
   679 => x"d40c8853",
   680 => x"bc905280",
   681 => x"c4d25193",
   682 => x"882d80c0",
   683 => x"e408762e",
   684 => x"09810689",
   685 => x"3880c0e4",
   686 => x"0880cad4",
   687 => x"0c8853bc",
   688 => x"9c5280c4",
   689 => x"ee519388",
   690 => x"2d80c0e4",
   691 => x"08893880",
   692 => x"c0e40880",
   693 => x"cad40c80",
   694 => x"cad40880",
   695 => x"2e818038",
   696 => x"80c7e20b",
   697 => x"80f52d80",
   698 => x"c7e30b80",
   699 => x"f52d7198",
   700 => x"2b71902b",
   701 => x"0780c7e4",
   702 => x"0b80f52d",
   703 => x"70882b72",
   704 => x"0780c7e5",
   705 => x"0b80f52d",
   706 => x"710780c8",
   707 => x"9a0b80f5",
   708 => x"2d80c89b",
   709 => x"0b80f52d",
   710 => x"71882b07",
   711 => x"535f5452",
   712 => x"5a565755",
   713 => x"7381abaa",
   714 => x"2e098106",
   715 => x"8e387551",
   716 => x"a9e22d80",
   717 => x"c0e40856",
   718 => x"96c80473",
   719 => x"82d4d52e",
   720 => x"8738bca8",
   721 => x"51979104",
   722 => x"80c49c52",
   723 => x"7551a8bf",
   724 => x"2d80c0e4",
   725 => x"085580c0",
   726 => x"e408802e",
   727 => x"83f73888",
   728 => x"53bc9c52",
   729 => x"80c4ee51",
   730 => x"93882d80",
   731 => x"c0e4088a",
   732 => x"38810b80",
   733 => x"caa80c97",
   734 => x"97048853",
   735 => x"bc905280",
   736 => x"c4d25193",
   737 => x"882d80c0",
   738 => x"e408802e",
   739 => x"8a38bcbc",
   740 => x"5186922d",
   741 => x"97f60480",
   742 => x"c89a0b80",
   743 => x"f52d5473",
   744 => x"80d52e09",
   745 => x"810680ce",
   746 => x"3880c89b",
   747 => x"0b80f52d",
   748 => x"547381aa",
   749 => x"2e098106",
   750 => x"bd38800b",
   751 => x"80c49c0b",
   752 => x"80f52d56",
   753 => x"547481e9",
   754 => x"2e833881",
   755 => x"547481eb",
   756 => x"2e8c3880",
   757 => x"5573752e",
   758 => x"09810682",
   759 => x"f83880c4",
   760 => x"a70b80f5",
   761 => x"2d55748e",
   762 => x"3880c4a8",
   763 => x"0b80f52d",
   764 => x"5473822e",
   765 => x"86388055",
   766 => x"9ad50480",
   767 => x"c4a90b80",
   768 => x"f52d7080",
   769 => x"caa00cff",
   770 => x"0580caa4",
   771 => x"0c80c4aa",
   772 => x"0b80f52d",
   773 => x"80c4ab0b",
   774 => x"80f52d58",
   775 => x"76057782",
   776 => x"80290570",
   777 => x"80cab00c",
   778 => x"80c4ac0b",
   779 => x"80f52d70",
   780 => x"80cac40c",
   781 => x"80caa808",
   782 => x"59575876",
   783 => x"802e81b6",
   784 => x"388853bc",
   785 => x"9c5280c4",
   786 => x"ee519388",
   787 => x"2d80c0e4",
   788 => x"08828238",
   789 => x"80caa008",
   790 => x"70842b80",
   791 => x"caac0c70",
   792 => x"80cac00c",
   793 => x"80c4c10b",
   794 => x"80f52d80",
   795 => x"c4c00b80",
   796 => x"f52d7182",
   797 => x"80290580",
   798 => x"c4c20b80",
   799 => x"f52d7084",
   800 => x"80802912",
   801 => x"80c4c30b",
   802 => x"80f52d70",
   803 => x"81800a29",
   804 => x"127080ca",
   805 => x"c80c80ca",
   806 => x"c4087129",
   807 => x"80cab008",
   808 => x"057080ca",
   809 => x"b40c80c4",
   810 => x"c90b80f5",
   811 => x"2d80c4c8",
   812 => x"0b80f52d",
   813 => x"71828029",
   814 => x"0580c4ca",
   815 => x"0b80f52d",
   816 => x"70848080",
   817 => x"291280c4",
   818 => x"cb0b80f5",
   819 => x"2d70982b",
   820 => x"81f00a06",
   821 => x"72057080",
   822 => x"cab80cfe",
   823 => x"117e2977",
   824 => x"0580cabc",
   825 => x"0c525952",
   826 => x"43545e51",
   827 => x"5259525d",
   828 => x"5759579a",
   829 => x"ce0480c4",
   830 => x"ae0b80f5",
   831 => x"2d80c4ad",
   832 => x"0b80f52d",
   833 => x"71828029",
   834 => x"057080ca",
   835 => x"ac0c70a0",
   836 => x"2983ff05",
   837 => x"70892a70",
   838 => x"80cac00c",
   839 => x"80c4b30b",
   840 => x"80f52d80",
   841 => x"c4b20b80",
   842 => x"f52d7182",
   843 => x"80290570",
   844 => x"80cac80c",
   845 => x"7b71291e",
   846 => x"7080cabc",
   847 => x"0c7d80ca",
   848 => x"b80c7305",
   849 => x"80cab40c",
   850 => x"555e5151",
   851 => x"55558051",
   852 => x"93c72d81",
   853 => x"557480c0",
   854 => x"e40c02a8",
   855 => x"050d0402",
   856 => x"ec050d76",
   857 => x"70872c71",
   858 => x"80ff0655",
   859 => x"565480ca",
   860 => x"a8088a38",
   861 => x"73882c74",
   862 => x"81ff0654",
   863 => x"5580c49c",
   864 => x"5280cab0",
   865 => x"081551a8",
   866 => x"bf2d80c0",
   867 => x"e4085480",
   868 => x"c0e40880",
   869 => x"2eb83880",
   870 => x"caa80880",
   871 => x"2e9a3872",
   872 => x"842980c4",
   873 => x"9c057008",
   874 => x"5253a9e2",
   875 => x"2d80c0e4",
   876 => x"08f00a06",
   877 => x"539bcc04",
   878 => x"721080c4",
   879 => x"9c057080",
   880 => x"e02d5253",
   881 => x"aa932d80",
   882 => x"c0e40853",
   883 => x"72547380",
   884 => x"c0e40c02",
   885 => x"94050d04",
   886 => x"02e0050d",
   887 => x"7970842c",
   888 => x"80cad008",
   889 => x"05718f06",
   890 => x"52555372",
   891 => x"8a3880c4",
   892 => x"9c527351",
   893 => x"a8bf2d72",
   894 => x"a02980c4",
   895 => x"9c055480",
   896 => x"7480f52d",
   897 => x"56537473",
   898 => x"2e833881",
   899 => x"537481e5",
   900 => x"2e81f438",
   901 => x"81707406",
   902 => x"54587280",
   903 => x"2e81e838",
   904 => x"8b1480f5",
   905 => x"2d70832a",
   906 => x"79065856",
   907 => x"769b3880",
   908 => x"c0940853",
   909 => x"72893872",
   910 => x"80c89c0b",
   911 => x"81b72d76",
   912 => x"80c0940c",
   913 => x"73539e89",
   914 => x"04758f2e",
   915 => x"09810681",
   916 => x"b638749f",
   917 => x"068d2980",
   918 => x"c88f1151",
   919 => x"53811480",
   920 => x"f52d7370",
   921 => x"81055581",
   922 => x"b72d8314",
   923 => x"80f52d73",
   924 => x"70810555",
   925 => x"81b72d85",
   926 => x"1480f52d",
   927 => x"73708105",
   928 => x"5581b72d",
   929 => x"871480f5",
   930 => x"2d737081",
   931 => x"055581b7",
   932 => x"2d891480",
   933 => x"f52d7370",
   934 => x"81055581",
   935 => x"b72d8e14",
   936 => x"80f52d73",
   937 => x"70810555",
   938 => x"81b72d90",
   939 => x"1480f52d",
   940 => x"73708105",
   941 => x"5581b72d",
   942 => x"921480f5",
   943 => x"2d737081",
   944 => x"055581b7",
   945 => x"2d941480",
   946 => x"f52d7370",
   947 => x"81055581",
   948 => x"b72d9614",
   949 => x"80f52d73",
   950 => x"70810555",
   951 => x"81b72d98",
   952 => x"1480f52d",
   953 => x"73708105",
   954 => x"5581b72d",
   955 => x"9c1480f5",
   956 => x"2d737081",
   957 => x"055581b7",
   958 => x"2d9e1480",
   959 => x"f52d7381",
   960 => x"b72d7780",
   961 => x"c0940c80",
   962 => x"537280c0",
   963 => x"e40c02a0",
   964 => x"050d0402",
   965 => x"cc050d7e",
   966 => x"605e5a80",
   967 => x"0b80cacc",
   968 => x"0880cad0",
   969 => x"08595c56",
   970 => x"805880ca",
   971 => x"ac08782e",
   972 => x"81b83877",
   973 => x"8f06a017",
   974 => x"57547391",
   975 => x"3880c49c",
   976 => x"52765181",
   977 => x"1757a8bf",
   978 => x"2d80c49c",
   979 => x"56807680",
   980 => x"f52d5654",
   981 => x"74742e83",
   982 => x"38815474",
   983 => x"81e52e80",
   984 => x"fd388170",
   985 => x"7506555c",
   986 => x"73802e80",
   987 => x"f1388b16",
   988 => x"80f52d98",
   989 => x"06597880",
   990 => x"e5388b53",
   991 => x"7c527551",
   992 => x"93882d80",
   993 => x"c0e40880",
   994 => x"d5389c16",
   995 => x"0851a9e2",
   996 => x"2d80c0e4",
   997 => x"08841b0c",
   998 => x"9a1680e0",
   999 => x"2d51aa93",
  1000 => x"2d80c0e4",
  1001 => x"0880c0e4",
  1002 => x"08881c0c",
  1003 => x"80c0e408",
  1004 => x"555580ca",
  1005 => x"a808802e",
  1006 => x"99389416",
  1007 => x"80e02d51",
  1008 => x"aa932d80",
  1009 => x"c0e40890",
  1010 => x"2b83fff0",
  1011 => x"0a067016",
  1012 => x"51547388",
  1013 => x"1b0c787a",
  1014 => x"0c7b54a0",
  1015 => x"a6048118",
  1016 => x"5880caac",
  1017 => x"087826fe",
  1018 => x"ca3880ca",
  1019 => x"a808802e",
  1020 => x"b3387a51",
  1021 => x"9adf2d80",
  1022 => x"c0e40880",
  1023 => x"c0e40880",
  1024 => x"fffffff8",
  1025 => x"06555b73",
  1026 => x"80ffffff",
  1027 => x"f82e9538",
  1028 => x"80c0e408",
  1029 => x"fe0580ca",
  1030 => x"a0082980",
  1031 => x"cab40805",
  1032 => x"579ea804",
  1033 => x"80547380",
  1034 => x"c0e40c02",
  1035 => x"b4050d04",
  1036 => x"02f4050d",
  1037 => x"74700881",
  1038 => x"05710c70",
  1039 => x"0880caa4",
  1040 => x"08065353",
  1041 => x"718f3888",
  1042 => x"1308519a",
  1043 => x"df2d80c0",
  1044 => x"e4088814",
  1045 => x"0c810b80",
  1046 => x"c0e40c02",
  1047 => x"8c050d04",
  1048 => x"02f0050d",
  1049 => x"75881108",
  1050 => x"fe0580ca",
  1051 => x"a0082980",
  1052 => x"cab40811",
  1053 => x"720880ca",
  1054 => x"a4080605",
  1055 => x"79555354",
  1056 => x"54a8bf2d",
  1057 => x"0290050d",
  1058 => x"0402f005",
  1059 => x"0d758811",
  1060 => x"08fe0580",
  1061 => x"caa00829",
  1062 => x"80cab408",
  1063 => x"11720880",
  1064 => x"caa40806",
  1065 => x"05795553",
  1066 => x"5454a6fd",
  1067 => x"2d029005",
  1068 => x"0d0402f4",
  1069 => x"050dd452",
  1070 => x"81ff720c",
  1071 => x"71085381",
  1072 => x"ff720c72",
  1073 => x"882b83fe",
  1074 => x"80067208",
  1075 => x"7081ff06",
  1076 => x"51525381",
  1077 => x"ff720c72",
  1078 => x"7107882b",
  1079 => x"72087081",
  1080 => x"ff065152",
  1081 => x"5381ff72",
  1082 => x"0c727107",
  1083 => x"882b7208",
  1084 => x"7081ff06",
  1085 => x"720780c0",
  1086 => x"e40c5253",
  1087 => x"028c050d",
  1088 => x"0402f405",
  1089 => x"0d747671",
  1090 => x"81ff06d4",
  1091 => x"0c535380",
  1092 => x"cad80885",
  1093 => x"3871892b",
  1094 => x"5271982a",
  1095 => x"d40c7190",
  1096 => x"2a7081ff",
  1097 => x"06d40c51",
  1098 => x"71882a70",
  1099 => x"81ff06d4",
  1100 => x"0c517181",
  1101 => x"ff06d40c",
  1102 => x"72902a70",
  1103 => x"81ff06d4",
  1104 => x"0c51d408",
  1105 => x"7081ff06",
  1106 => x"515182b8",
  1107 => x"bf527081",
  1108 => x"ff2e0981",
  1109 => x"06943881",
  1110 => x"ff0bd40c",
  1111 => x"d4087081",
  1112 => x"ff06ff14",
  1113 => x"54515171",
  1114 => x"e5387080",
  1115 => x"c0e40c02",
  1116 => x"8c050d04",
  1117 => x"02fc050d",
  1118 => x"81c75181",
  1119 => x"ff0bd40c",
  1120 => x"ff115170",
  1121 => x"8025f438",
  1122 => x"0284050d",
  1123 => x"0402f005",
  1124 => x"0da2f42d",
  1125 => x"8fcf5380",
  1126 => x"5287fc80",
  1127 => x"f751a281",
  1128 => x"2d80c0e4",
  1129 => x"085480c0",
  1130 => x"e408812e",
  1131 => x"098106a4",
  1132 => x"3881ff0b",
  1133 => x"d40c820a",
  1134 => x"52849c80",
  1135 => x"e951a281",
  1136 => x"2d80c0e4",
  1137 => x"088b3881",
  1138 => x"ff0bd40c",
  1139 => x"7353a3db",
  1140 => x"04a2f42d",
  1141 => x"ff135372",
  1142 => x"ffbd3872",
  1143 => x"80c0e40c",
  1144 => x"0290050d",
  1145 => x"0402f405",
  1146 => x"0d81ff0b",
  1147 => x"d40c9353",
  1148 => x"805287fc",
  1149 => x"80c151a2",
  1150 => x"812d80c0",
  1151 => x"e4088b38",
  1152 => x"81ff0bd4",
  1153 => x"0c8153a4",
  1154 => x"9304a2f4",
  1155 => x"2dff1353",
  1156 => x"72de3872",
  1157 => x"80c0e40c",
  1158 => x"028c050d",
  1159 => x"0402f005",
  1160 => x"0da2f42d",
  1161 => x"83aa5284",
  1162 => x"9c80c851",
  1163 => x"a2812d80",
  1164 => x"c0e40881",
  1165 => x"2e098106",
  1166 => x"9338a1b2",
  1167 => x"2d80c0e4",
  1168 => x"0883ffff",
  1169 => x"06537283",
  1170 => x"aa2e9738",
  1171 => x"a3e52da4",
  1172 => x"dd048154",
  1173 => x"a5c504bc",
  1174 => x"c8518692",
  1175 => x"2d8054a5",
  1176 => x"c50481ff",
  1177 => x"0bd40cb1",
  1178 => x"53a38d2d",
  1179 => x"80c0e408",
  1180 => x"802e80c2",
  1181 => x"38805287",
  1182 => x"fc80fa51",
  1183 => x"a2812d80",
  1184 => x"c0e408b2",
  1185 => x"3881ff0b",
  1186 => x"d40cd408",
  1187 => x"5381ff0b",
  1188 => x"d40c81ff",
  1189 => x"0bd40c81",
  1190 => x"ff0bd40c",
  1191 => x"81ff0bd4",
  1192 => x"0c72862a",
  1193 => x"70810680",
  1194 => x"c0e40856",
  1195 => x"51537280",
  1196 => x"2e9338a4",
  1197 => x"d2047282",
  1198 => x"2eff9c38",
  1199 => x"ff135372",
  1200 => x"ffa73872",
  1201 => x"547380c0",
  1202 => x"e40c0290",
  1203 => x"050d0402",
  1204 => x"f0050d81",
  1205 => x"0b80cad8",
  1206 => x"0c8454d0",
  1207 => x"08708f2a",
  1208 => x"70810651",
  1209 => x"515372f3",
  1210 => x"3872d00c",
  1211 => x"a2f42dbc",
  1212 => x"d8518692",
  1213 => x"2dd00870",
  1214 => x"8f2a7081",
  1215 => x"06515153",
  1216 => x"72f33881",
  1217 => x"0bd00cb1",
  1218 => x"53805284",
  1219 => x"d480c051",
  1220 => x"a2812d80",
  1221 => x"c0e40881",
  1222 => x"2ea13872",
  1223 => x"822e0981",
  1224 => x"068c38bc",
  1225 => x"e4518692",
  1226 => x"2d8053a6",
  1227 => x"f304ff13",
  1228 => x"5372d638",
  1229 => x"ff145473",
  1230 => x"ffa138a4",
  1231 => x"9d2d80c0",
  1232 => x"e40880ca",
  1233 => x"d80c80c0",
  1234 => x"e4088b38",
  1235 => x"815287fc",
  1236 => x"80d051a2",
  1237 => x"812d81ff",
  1238 => x"0bd40cd0",
  1239 => x"08708f2a",
  1240 => x"70810651",
  1241 => x"515372f3",
  1242 => x"3872d00c",
  1243 => x"81ff0bd4",
  1244 => x"0c815372",
  1245 => x"80c0e40c",
  1246 => x"0290050d",
  1247 => x"0402e805",
  1248 => x"0d785681",
  1249 => x"ff0bd40c",
  1250 => x"d008708f",
  1251 => x"2a708106",
  1252 => x"51515372",
  1253 => x"f3388281",
  1254 => x"0bd00c81",
  1255 => x"ff0bd40c",
  1256 => x"775287fc",
  1257 => x"80d851a2",
  1258 => x"812d80c0",
  1259 => x"e408802e",
  1260 => x"8c38bcfc",
  1261 => x"5186922d",
  1262 => x"8153a8b5",
  1263 => x"0481ff0b",
  1264 => x"d40c81fe",
  1265 => x"0bd40c80",
  1266 => x"ff557570",
  1267 => x"84055708",
  1268 => x"70982ad4",
  1269 => x"0c70902c",
  1270 => x"7081ff06",
  1271 => x"d40c5470",
  1272 => x"882c7081",
  1273 => x"ff06d40c",
  1274 => x"547081ff",
  1275 => x"06d40c54",
  1276 => x"ff155574",
  1277 => x"8025d338",
  1278 => x"81ff0bd4",
  1279 => x"0c81ff0b",
  1280 => x"d40c81ff",
  1281 => x"0bd40c86",
  1282 => x"8da05481",
  1283 => x"ff0bd40c",
  1284 => x"d40881ff",
  1285 => x"06557487",
  1286 => x"38ff1454",
  1287 => x"73ed3881",
  1288 => x"ff0bd40c",
  1289 => x"d008708f",
  1290 => x"2a708106",
  1291 => x"51515372",
  1292 => x"f33872d0",
  1293 => x"0c7280c0",
  1294 => x"e40c0298",
  1295 => x"050d0402",
  1296 => x"e8050d78",
  1297 => x"55805681",
  1298 => x"ff0bd40c",
  1299 => x"d008708f",
  1300 => x"2a708106",
  1301 => x"51515372",
  1302 => x"f3388281",
  1303 => x"0bd00c81",
  1304 => x"ff0bd40c",
  1305 => x"775287fc",
  1306 => x"80d151a2",
  1307 => x"812d80db",
  1308 => x"c6df5480",
  1309 => x"c0e40880",
  1310 => x"2e8a38bd",
  1311 => x"8c518692",
  1312 => x"2da9d804",
  1313 => x"81ff0bd4",
  1314 => x"0cd40870",
  1315 => x"81ff0651",
  1316 => x"537281fe",
  1317 => x"2e098106",
  1318 => x"9e3880ff",
  1319 => x"53a1b22d",
  1320 => x"80c0e408",
  1321 => x"75708405",
  1322 => x"570cff13",
  1323 => x"53728025",
  1324 => x"ec388156",
  1325 => x"a9bd04ff",
  1326 => x"145473c8",
  1327 => x"3881ff0b",
  1328 => x"d40c81ff",
  1329 => x"0bd40cd0",
  1330 => x"08708f2a",
  1331 => x"70810651",
  1332 => x"515372f3",
  1333 => x"3872d00c",
  1334 => x"7580c0e4",
  1335 => x"0c029805",
  1336 => x"0d0402f4",
  1337 => x"050d7470",
  1338 => x"882a83fe",
  1339 => x"80067072",
  1340 => x"982a0772",
  1341 => x"882b87fc",
  1342 => x"80800673",
  1343 => x"982b81f0",
  1344 => x"0a067173",
  1345 => x"070780c0",
  1346 => x"e40c5651",
  1347 => x"5351028c",
  1348 => x"050d0402",
  1349 => x"f8050d02",
  1350 => x"8e0580f5",
  1351 => x"2d74882b",
  1352 => x"077083ff",
  1353 => x"ff0680c0",
  1354 => x"e40c5102",
  1355 => x"88050d04",
  1356 => x"02fc050d",
  1357 => x"72518071",
  1358 => x"0c800b84",
  1359 => x"120c0284",
  1360 => x"050d0402",
  1361 => x"f0050d75",
  1362 => x"70088412",
  1363 => x"08535353",
  1364 => x"ff547171",
  1365 => x"2ea838ae",
  1366 => x"9a2d8413",
  1367 => x"08708429",
  1368 => x"14881170",
  1369 => x"087081ff",
  1370 => x"06841808",
  1371 => x"81118706",
  1372 => x"841a0c53",
  1373 => x"51555151",
  1374 => x"51ae942d",
  1375 => x"71547380",
  1376 => x"c0e40c02",
  1377 => x"90050d04",
  1378 => x"02f8050d",
  1379 => x"ae9a2de0",
  1380 => x"08708b2a",
  1381 => x"70810651",
  1382 => x"52527080",
  1383 => x"2ea13880",
  1384 => x"cadc0870",
  1385 => x"842980ca",
  1386 => x"e4057381",
  1387 => x"ff06710c",
  1388 => x"515180ca",
  1389 => x"dc088111",
  1390 => x"870680ca",
  1391 => x"dc0c5180",
  1392 => x"0b80cb84",
  1393 => x"0cae8c2d",
  1394 => x"ae942d02",
  1395 => x"88050d04",
  1396 => x"02fc050d",
  1397 => x"ae9a2d81",
  1398 => x"0b80cb84",
  1399 => x"0cae942d",
  1400 => x"80cb8408",
  1401 => x"5170f938",
  1402 => x"0284050d",
  1403 => x"0402fc05",
  1404 => x"0d80cadc",
  1405 => x"51aab02d",
  1406 => x"ab8851ae",
  1407 => x"882dadaf",
  1408 => x"2d028405",
  1409 => x"0d0402f4",
  1410 => x"050dad94",
  1411 => x"0480c0e4",
  1412 => x"0881f02e",
  1413 => x"0981068a",
  1414 => x"38810b80",
  1415 => x"c0d80cad",
  1416 => x"940480c0",
  1417 => x"e40881e0",
  1418 => x"2e098106",
  1419 => x"8a38810b",
  1420 => x"80c0dc0c",
  1421 => x"ad940480",
  1422 => x"c0e40852",
  1423 => x"80c0dc08",
  1424 => x"802e8938",
  1425 => x"80c0e408",
  1426 => x"81800552",
  1427 => x"71842c72",
  1428 => x"8f065353",
  1429 => x"80c0d808",
  1430 => x"802e9a38",
  1431 => x"72842980",
  1432 => x"c0980572",
  1433 => x"1381712b",
  1434 => x"70097308",
  1435 => x"06730c51",
  1436 => x"5353ad88",
  1437 => x"04728429",
  1438 => x"80c09805",
  1439 => x"72138371",
  1440 => x"2b720807",
  1441 => x"720c5353",
  1442 => x"800b80c0",
  1443 => x"dc0c800b",
  1444 => x"80c0d80c",
  1445 => x"80cadc51",
  1446 => x"aac32d80",
  1447 => x"c0e408ff",
  1448 => x"24feea38",
  1449 => x"800b80c0",
  1450 => x"e40c028c",
  1451 => x"050d0402",
  1452 => x"f8050d80",
  1453 => x"c098528f",
  1454 => x"51807270",
  1455 => x"8405540c",
  1456 => x"ff115170",
  1457 => x"8025f238",
  1458 => x"0288050d",
  1459 => x"0402f005",
  1460 => x"0d7551ae",
  1461 => x"9a2d7082",
  1462 => x"2cfc0680",
  1463 => x"c0981172",
  1464 => x"109e0671",
  1465 => x"0870722a",
  1466 => x"70830682",
  1467 => x"742b7009",
  1468 => x"7406760c",
  1469 => x"54515657",
  1470 => x"535153ae",
  1471 => x"942d7180",
  1472 => x"c0e40c02",
  1473 => x"90050d04",
  1474 => x"71980c04",
  1475 => x"ffb00880",
  1476 => x"c0e40c04",
  1477 => x"810bffb0",
  1478 => x"0c04800b",
  1479 => x"ffb00c04",
  1480 => x"02fc050d",
  1481 => x"810b80c0",
  1482 => x"e00c8151",
  1483 => x"85812d02",
  1484 => x"84050d04",
  1485 => x"02fc050d",
  1486 => x"800b80c0",
  1487 => x"e00c8051",
  1488 => x"85812d02",
  1489 => x"84050d04",
  1490 => x"02ec050d",
  1491 => x"76548052",
  1492 => x"870b8815",
  1493 => x"80f52d56",
  1494 => x"53747224",
  1495 => x"8338a053",
  1496 => x"725182f8",
  1497 => x"2d81128b",
  1498 => x"1580f52d",
  1499 => x"54527272",
  1500 => x"25de3802",
  1501 => x"94050d04",
  1502 => x"02f0050d",
  1503 => x"80cb9408",
  1504 => x"5481f92d",
  1505 => x"800b80cb",
  1506 => x"980c7308",
  1507 => x"802e8186",
  1508 => x"38820b80",
  1509 => x"c0f80c80",
  1510 => x"cb98088f",
  1511 => x"0680c0f4",
  1512 => x"0c730852",
  1513 => x"71832e96",
  1514 => x"38718326",
  1515 => x"89387181",
  1516 => x"2eaf38af",
  1517 => x"ff047185",
  1518 => x"2e9f38af",
  1519 => x"ff048814",
  1520 => x"80f52d84",
  1521 => x"1508bd9c",
  1522 => x"53545286",
  1523 => x"922d7184",
  1524 => x"29137008",
  1525 => x"5252b083",
  1526 => x"047351ae",
  1527 => x"c82dafff",
  1528 => x"0480cb88",
  1529 => x"08881508",
  1530 => x"2c708106",
  1531 => x"51527180",
  1532 => x"2e8738bd",
  1533 => x"a051affc",
  1534 => x"04bda451",
  1535 => x"86922d84",
  1536 => x"14085186",
  1537 => x"922d80cb",
  1538 => x"98088105",
  1539 => x"80cb980c",
  1540 => x"8c1454af",
  1541 => x"8a040290",
  1542 => x"050d0471",
  1543 => x"80cb940c",
  1544 => x"aef82d80",
  1545 => x"cb9808ff",
  1546 => x"0580cb9c",
  1547 => x"0c0402e8",
  1548 => x"050d80cb",
  1549 => x"940880cb",
  1550 => x"a0085755",
  1551 => x"80f851ad",
  1552 => x"cd2d80c0",
  1553 => x"e408812a",
  1554 => x"70810651",
  1555 => x"52719c38",
  1556 => x"8751adcd",
  1557 => x"2d80c0e4",
  1558 => x"08812a70",
  1559 => x"81065152",
  1560 => x"71802eb5",
  1561 => x"38b0eb04",
  1562 => x"ac862d87",
  1563 => x"51adcd2d",
  1564 => x"80c0e408",
  1565 => x"f338b0fc",
  1566 => x"04ac862d",
  1567 => x"80f851ad",
  1568 => x"cd2d80c0",
  1569 => x"e408f238",
  1570 => x"80c0e008",
  1571 => x"81327080",
  1572 => x"c0e00c70",
  1573 => x"52528581",
  1574 => x"2d800b80",
  1575 => x"cb8c0c80",
  1576 => x"0b80cb90",
  1577 => x"0c80c0e0",
  1578 => x"08838d38",
  1579 => x"80da51ad",
  1580 => x"cd2d80c0",
  1581 => x"e408802e",
  1582 => x"8c3880cb",
  1583 => x"8c088180",
  1584 => x"0780cb8c",
  1585 => x"0c80d951",
  1586 => x"adcd2d80",
  1587 => x"c0e40880",
  1588 => x"2e8c3880",
  1589 => x"cb8c0880",
  1590 => x"c00780cb",
  1591 => x"8c0c8194",
  1592 => x"51adcd2d",
  1593 => x"80c0e408",
  1594 => x"802e8b38",
  1595 => x"80cb8c08",
  1596 => x"900780cb",
  1597 => x"8c0c8191",
  1598 => x"51adcd2d",
  1599 => x"80c0e408",
  1600 => x"802e8b38",
  1601 => x"80cb8c08",
  1602 => x"a00780cb",
  1603 => x"8c0c81f5",
  1604 => x"51adcd2d",
  1605 => x"80c0e408",
  1606 => x"802e8b38",
  1607 => x"80cb8c08",
  1608 => x"810780cb",
  1609 => x"8c0c81f2",
  1610 => x"51adcd2d",
  1611 => x"80c0e408",
  1612 => x"802e8b38",
  1613 => x"80cb8c08",
  1614 => x"820780cb",
  1615 => x"8c0c81eb",
  1616 => x"51adcd2d",
  1617 => x"80c0e408",
  1618 => x"802e8b38",
  1619 => x"80cb8c08",
  1620 => x"840780cb",
  1621 => x"8c0c81f4",
  1622 => x"51adcd2d",
  1623 => x"80c0e408",
  1624 => x"802e8b38",
  1625 => x"80cb8c08",
  1626 => x"880780cb",
  1627 => x"8c0c80d8",
  1628 => x"51adcd2d",
  1629 => x"80c0e408",
  1630 => x"802e8c38",
  1631 => x"80cb9008",
  1632 => x"81800780",
  1633 => x"cb900c92",
  1634 => x"51adcd2d",
  1635 => x"80c0e408",
  1636 => x"802e8c38",
  1637 => x"80cb9008",
  1638 => x"80c00780",
  1639 => x"cb900c94",
  1640 => x"51adcd2d",
  1641 => x"80c0e408",
  1642 => x"802e8b38",
  1643 => x"80cb9008",
  1644 => x"900780cb",
  1645 => x"900c9151",
  1646 => x"adcd2d80",
  1647 => x"c0e40880",
  1648 => x"2e8b3880",
  1649 => x"cb9008a0",
  1650 => x"0780cb90",
  1651 => x"0c9d51ad",
  1652 => x"cd2d80c0",
  1653 => x"e408802e",
  1654 => x"8b3880cb",
  1655 => x"90088107",
  1656 => x"80cb900c",
  1657 => x"9b51adcd",
  1658 => x"2d80c0e4",
  1659 => x"08802e8b",
  1660 => x"3880cb90",
  1661 => x"08820780",
  1662 => x"cb900c9c",
  1663 => x"51adcd2d",
  1664 => x"80c0e408",
  1665 => x"802e8b38",
  1666 => x"80cb9008",
  1667 => x"840780cb",
  1668 => x"900ca351",
  1669 => x"adcd2d80",
  1670 => x"c0e40880",
  1671 => x"2e8b3880",
  1672 => x"cb900888",
  1673 => x"0780cb90",
  1674 => x"0c81fd51",
  1675 => x"adcd2d81",
  1676 => x"fa51adcd",
  1677 => x"2dba8d04",
  1678 => x"81f551ad",
  1679 => x"cd2d80c0",
  1680 => x"e408812a",
  1681 => x"70810651",
  1682 => x"5271802e",
  1683 => x"b33880cb",
  1684 => x"9c085271",
  1685 => x"802e8a38",
  1686 => x"ff1280cb",
  1687 => x"9c0cb580",
  1688 => x"0480cb98",
  1689 => x"081080cb",
  1690 => x"98080570",
  1691 => x"84291651",
  1692 => x"52881208",
  1693 => x"802e8938",
  1694 => x"ff518812",
  1695 => x"0852712d",
  1696 => x"81f251ad",
  1697 => x"cd2d80c0",
  1698 => x"e408812a",
  1699 => x"70810651",
  1700 => x"5271802e",
  1701 => x"b43880cb",
  1702 => x"9808ff11",
  1703 => x"80cb9c08",
  1704 => x"56535373",
  1705 => x"72258a38",
  1706 => x"811480cb",
  1707 => x"9c0cb5c9",
  1708 => x"04721013",
  1709 => x"70842916",
  1710 => x"51528812",
  1711 => x"08802e89",
  1712 => x"38fe5188",
  1713 => x"12085271",
  1714 => x"2d81fd51",
  1715 => x"adcd2d80",
  1716 => x"c0e40881",
  1717 => x"2a708106",
  1718 => x"51527180",
  1719 => x"2eb13880",
  1720 => x"cb9c0880",
  1721 => x"2e8a3880",
  1722 => x"0b80cb9c",
  1723 => x"0cb68f04",
  1724 => x"80cb9808",
  1725 => x"1080cb98",
  1726 => x"08057084",
  1727 => x"29165152",
  1728 => x"88120880",
  1729 => x"2e8938fd",
  1730 => x"51881208",
  1731 => x"52712d81",
  1732 => x"fa51adcd",
  1733 => x"2d80c0e4",
  1734 => x"08812a70",
  1735 => x"81065152",
  1736 => x"71802eb1",
  1737 => x"3880cb98",
  1738 => x"08ff1154",
  1739 => x"5280cb9c",
  1740 => x"08732589",
  1741 => x"387280cb",
  1742 => x"9c0cb6d5",
  1743 => x"04711012",
  1744 => x"70842916",
  1745 => x"51528812",
  1746 => x"08802e89",
  1747 => x"38fc5188",
  1748 => x"12085271",
  1749 => x"2d80cb9c",
  1750 => x"08705354",
  1751 => x"73802e8a",
  1752 => x"388c15ff",
  1753 => x"155555b6",
  1754 => x"dc04820b",
  1755 => x"80c0f80c",
  1756 => x"718f0680",
  1757 => x"c0f40c81",
  1758 => x"eb51adcd",
  1759 => x"2d80c0e4",
  1760 => x"08812a70",
  1761 => x"81065152",
  1762 => x"71802ead",
  1763 => x"38740885",
  1764 => x"2e098106",
  1765 => x"a4388815",
  1766 => x"80f52dff",
  1767 => x"05527188",
  1768 => x"1681b72d",
  1769 => x"71982b52",
  1770 => x"71802588",
  1771 => x"38800b88",
  1772 => x"1681b72d",
  1773 => x"7451aec8",
  1774 => x"2d81f451",
  1775 => x"adcd2d80",
  1776 => x"c0e40881",
  1777 => x"2a708106",
  1778 => x"51527180",
  1779 => x"2eb33874",
  1780 => x"08852e09",
  1781 => x"8106aa38",
  1782 => x"881580f5",
  1783 => x"2d810552",
  1784 => x"71881681",
  1785 => x"b72d7181",
  1786 => x"ff068b16",
  1787 => x"80f52d54",
  1788 => x"52727227",
  1789 => x"87387288",
  1790 => x"1681b72d",
  1791 => x"7451aec8",
  1792 => x"2d80da51",
  1793 => x"adcd2d80",
  1794 => x"c0e40881",
  1795 => x"2a708106",
  1796 => x"51527180",
  1797 => x"2e81ad38",
  1798 => x"80cb9408",
  1799 => x"80cb9c08",
  1800 => x"55537380",
  1801 => x"2e8a388c",
  1802 => x"13ff1555",
  1803 => x"53b8a204",
  1804 => x"72085271",
  1805 => x"822ea638",
  1806 => x"71822689",
  1807 => x"3871812e",
  1808 => x"aa38b9c4",
  1809 => x"0471832e",
  1810 => x"b4387184",
  1811 => x"2e098106",
  1812 => x"80f23888",
  1813 => x"130851b0",
  1814 => x"9b2db9c4",
  1815 => x"0480cb9c",
  1816 => x"08518813",
  1817 => x"0852712d",
  1818 => x"b9c40481",
  1819 => x"0b881408",
  1820 => x"2b80cb88",
  1821 => x"083280cb",
  1822 => x"880cb998",
  1823 => x"04881380",
  1824 => x"f52d8105",
  1825 => x"8b1480f5",
  1826 => x"2d535471",
  1827 => x"74248338",
  1828 => x"80547388",
  1829 => x"1481b72d",
  1830 => x"aef82db9",
  1831 => x"c4047508",
  1832 => x"802ea438",
  1833 => x"750851ad",
  1834 => x"cd2d80c0",
  1835 => x"e4088106",
  1836 => x"5271802e",
  1837 => x"8c3880cb",
  1838 => x"9c085184",
  1839 => x"16085271",
  1840 => x"2d881656",
  1841 => x"75d83880",
  1842 => x"54800b80",
  1843 => x"c0f80c73",
  1844 => x"8f0680c0",
  1845 => x"f40ca052",
  1846 => x"7380cb9c",
  1847 => x"082e0981",
  1848 => x"06993880",
  1849 => x"cb9808ff",
  1850 => x"05743270",
  1851 => x"09810570",
  1852 => x"72079f2a",
  1853 => x"91713151",
  1854 => x"51535371",
  1855 => x"5182f82d",
  1856 => x"8114548e",
  1857 => x"7425c238",
  1858 => x"80c0e008",
  1859 => x"527180c0",
  1860 => x"e40c0298",
  1861 => x"050d0400",
  1862 => x"00ffffff",
  1863 => x"ff00ffff",
  1864 => x"ffff00ff",
  1865 => x"ffffff00",
  1866 => x"4f4b0000",
  1867 => x"52657365",
  1868 => x"74000000",
  1869 => x"53617665",
  1870 => x"20736574",
  1871 => x"74696e67",
  1872 => x"73000000",
  1873 => x"5363616e",
  1874 => x"6c696e65",
  1875 => x"73000000",
  1876 => x"41756469",
  1877 => x"6f20566f",
  1878 => x"6c756d65",
  1879 => x"00000000",
  1880 => x"4c6f6164",
  1881 => x"20524f4d",
  1882 => x"20100000",
  1883 => x"45786974",
  1884 => x"00000000",
  1885 => x"4a6f7973",
  1886 => x"7469636b",
  1887 => x"20737761",
  1888 => x"70000000",
  1889 => x"4a6f7973",
  1890 => x"7469636b",
  1891 => x"206e6f72",
  1892 => x"6d616c00",
  1893 => x"56474120",
  1894 => x"2d203331",
  1895 => x"4b487a00",
  1896 => x"5456202d",
  1897 => x"2031354b",
  1898 => x"487a0000",
  1899 => x"4261636b",
  1900 => x"00000000",
  1901 => x"4c6f6164",
  1902 => x"20457272",
  1903 => x"6f722100",
  1904 => x"46504741",
  1905 => x"47454e20",
  1906 => x"43464700",
  1907 => x"496e6974",
  1908 => x"69616c69",
  1909 => x"7a696e67",
  1910 => x"20534420",
  1911 => x"63617264",
  1912 => x"0a000000",
  1913 => x"424f4f54",
  1914 => x"20202020",
  1915 => x"47454e00",
  1916 => x"43617264",
  1917 => x"20696e69",
  1918 => x"74206661",
  1919 => x"696c6564",
  1920 => x"0a000000",
  1921 => x"4d425220",
  1922 => x"6661696c",
  1923 => x"0a000000",
  1924 => x"46415431",
  1925 => x"36202020",
  1926 => x"00000000",
  1927 => x"46415433",
  1928 => x"32202020",
  1929 => x"00000000",
  1930 => x"4e6f2070",
  1931 => x"61727469",
  1932 => x"74696f6e",
  1933 => x"20736967",
  1934 => x"0a000000",
  1935 => x"42616420",
  1936 => x"70617274",
  1937 => x"0a000000",
  1938 => x"53444843",
  1939 => x"20657272",
  1940 => x"6f72210a",
  1941 => x"00000000",
  1942 => x"53442069",
  1943 => x"6e69742e",
  1944 => x"2e2e0a00",
  1945 => x"53442063",
  1946 => x"61726420",
  1947 => x"72657365",
  1948 => x"74206661",
  1949 => x"696c6564",
  1950 => x"210a0000",
  1951 => x"57726974",
  1952 => x"65206661",
  1953 => x"696c6564",
  1954 => x"0a000000",
  1955 => x"52656164",
  1956 => x"20666169",
  1957 => x"6c65640a",
  1958 => x"00000000",
  1959 => x"16200000",
  1960 => x"14200000",
  1961 => x"15200000",
  1962 => x"00000002",
  1963 => x"00000000",
  1964 => x"00000002",
  1965 => x"00001d2c",
  1966 => x"000004dd",
  1967 => x"00000002",
  1968 => x"00001d34",
  1969 => x"000003a2",
  1970 => x"00000003",
  1971 => x"00001f24",
  1972 => x"00000002",
  1973 => x"00000001",
  1974 => x"00001d44",
  1975 => x"00000001",
  1976 => x"00000003",
  1977 => x"00001f1c",
  1978 => x"00000002",
  1979 => x"00000005",
  1980 => x"00001d50",
  1981 => x"00000007",
  1982 => x"00000002",
  1983 => x"00001d60",
  1984 => x"000007a1",
  1985 => x"00000002",
  1986 => x"00001d6c",
  1987 => x"00001734",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000000",
  1991 => x"00001d74",
  1992 => x"00001d84",
  1993 => x"00001d94",
  1994 => x"00001da0",
  1995 => x"00000002",
  1996 => x"00002094",
  1997 => x"0000056f",
  1998 => x"00000002",
  1999 => x"000020b2",
  2000 => x"0000056f",
  2001 => x"00000002",
  2002 => x"000020d0",
  2003 => x"0000056f",
  2004 => x"00000002",
  2005 => x"000020ee",
  2006 => x"0000056f",
  2007 => x"00000002",
  2008 => x"0000210c",
  2009 => x"0000056f",
  2010 => x"00000002",
  2011 => x"0000212a",
  2012 => x"0000056f",
  2013 => x"00000002",
  2014 => x"00002148",
  2015 => x"0000056f",
  2016 => x"00000002",
  2017 => x"00002166",
  2018 => x"0000056f",
  2019 => x"00000002",
  2020 => x"00002184",
  2021 => x"0000056f",
  2022 => x"00000002",
  2023 => x"000021a2",
  2024 => x"0000056f",
  2025 => x"00000002",
  2026 => x"000021c0",
  2027 => x"0000056f",
  2028 => x"00000002",
  2029 => x"000021de",
  2030 => x"0000056f",
  2031 => x"00000002",
  2032 => x"000021fc",
  2033 => x"0000056f",
  2034 => x"00000004",
  2035 => x"00001dac",
  2036 => x"00001eb0",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000735",
  2040 => x"00000000",
  2041 => x"00000004",
  2042 => x"00001db4",
  2043 => x"00001eb0",
  2044 => x"00000004",
  2045 => x"00001e54",
  2046 => x"00001eb0",
  2047 => x"00000004",
  2048 => x"00001d28",
  2049 => x"00001eb0",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

